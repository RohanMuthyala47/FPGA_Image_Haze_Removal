module Transmission_Reciprocal_LUT (
    input      [13:0] in,  // Q0.14 input (unsigned, ranges from 0 to 0.65)
    output reg [11:0] out  // Q2.10 reciprocal output (unsigned, 12-bit)
);

    always @(*) begin
        case(in)
            14'd    0: out = 12'h400;
            14'd    1: out = 12'h400;
            14'd    2: out = 12'h400;
            14'd    3: out = 12'h400;
            14'd    4: out = 12'h400;
            14'd    5: out = 12'h400;
            14'd    6: out = 12'h400;
            14'd    7: out = 12'h400;
            14'd    8: out = 12'h401;
            14'd    9: out = 12'h401;
            14'd   10: out = 12'h401;
            14'd   11: out = 12'h401;
            14'd   12: out = 12'h401;
            14'd   13: out = 12'h401;
            14'd   14: out = 12'h401;
            14'd   15: out = 12'h401;
            14'd   16: out = 12'h401;
            14'd   17: out = 12'h401;
            14'd   18: out = 12'h401;
            14'd   19: out = 12'h401;
            14'd   20: out = 12'h401;
            14'd   21: out = 12'h401;
            14'd   22: out = 12'h401;
            14'd   23: out = 12'h401;
            14'd   24: out = 12'h402;
            14'd   25: out = 12'h402;
            14'd   26: out = 12'h402;
            14'd   27: out = 12'h402;
            14'd   28: out = 12'h402;
            14'd   29: out = 12'h402;
            14'd   30: out = 12'h402;
            14'd   31: out = 12'h402;
            14'd   32: out = 12'h402;
            14'd   33: out = 12'h402;
            14'd   34: out = 12'h402;
            14'd   35: out = 12'h402;
            14'd   36: out = 12'h402;
            14'd   37: out = 12'h402;
            14'd   38: out = 12'h402;
            14'd   39: out = 12'h402;
            14'd   40: out = 12'h403;
            14'd   41: out = 12'h403;
            14'd   42: out = 12'h403;
            14'd   43: out = 12'h403;
            14'd   44: out = 12'h403;
            14'd   45: out = 12'h403;
            14'd   46: out = 12'h403;
            14'd   47: out = 12'h403;
            14'd   48: out = 12'h403;
            14'd   49: out = 12'h403;
            14'd   50: out = 12'h403;
            14'd   51: out = 12'h403;
            14'd   52: out = 12'h403;
            14'd   53: out = 12'h403;
            14'd   54: out = 12'h403;
            14'd   55: out = 12'h403;
            14'd   56: out = 12'h404;
            14'd   57: out = 12'h404;
            14'd   58: out = 12'h404;
            14'd   59: out = 12'h404;
            14'd   60: out = 12'h404;
            14'd   61: out = 12'h404;
            14'd   62: out = 12'h404;
            14'd   63: out = 12'h404;
            14'd   64: out = 12'h404;
            14'd   65: out = 12'h404;
            14'd   66: out = 12'h404;
            14'd   67: out = 12'h404;
            14'd   68: out = 12'h404;
            14'd   69: out = 12'h404;
            14'd   70: out = 12'h404;
            14'd   71: out = 12'h404;
            14'd   72: out = 12'h405;
            14'd   73: out = 12'h405;
            14'd   74: out = 12'h405;
            14'd   75: out = 12'h405;
            14'd   76: out = 12'h405;
            14'd   77: out = 12'h405;
            14'd   78: out = 12'h405;
            14'd   79: out = 12'h405;
            14'd   80: out = 12'h405;
            14'd   81: out = 12'h405;
            14'd   82: out = 12'h405;
            14'd   83: out = 12'h405;
            14'd   84: out = 12'h405;
            14'd   85: out = 12'h405;
            14'd   86: out = 12'h405;
            14'd   87: out = 12'h405;
            14'd   88: out = 12'h406;
            14'd   89: out = 12'h406;
            14'd   90: out = 12'h406;
            14'd   91: out = 12'h406;
            14'd   92: out = 12'h406;
            14'd   93: out = 12'h406;
            14'd   94: out = 12'h406;
            14'd   95: out = 12'h406;
            14'd   96: out = 12'h406;
            14'd   97: out = 12'h406;
            14'd   98: out = 12'h406;
            14'd   99: out = 12'h406;
            14'd  100: out = 12'h406;
            14'd  101: out = 12'h406;
            14'd  102: out = 12'h406;
            14'd  103: out = 12'h406;
            14'd  104: out = 12'h407;
            14'd  105: out = 12'h407;
            14'd  106: out = 12'h407;
            14'd  107: out = 12'h407;
            14'd  108: out = 12'h407;
            14'd  109: out = 12'h407;
            14'd  110: out = 12'h407;
            14'd  111: out = 12'h407;
            14'd  112: out = 12'h407;
            14'd  113: out = 12'h407;
            14'd  114: out = 12'h407;
            14'd  115: out = 12'h407;
            14'd  116: out = 12'h407;
            14'd  117: out = 12'h407;
            14'd  118: out = 12'h407;
            14'd  119: out = 12'h407;
            14'd  120: out = 12'h408;
            14'd  121: out = 12'h408;
            14'd  122: out = 12'h408;
            14'd  123: out = 12'h408;
            14'd  124: out = 12'h408;
            14'd  125: out = 12'h408;
            14'd  126: out = 12'h408;
            14'd  127: out = 12'h408;
            14'd  128: out = 12'h408;
            14'd  129: out = 12'h408;
            14'd  130: out = 12'h408;
            14'd  131: out = 12'h408;
            14'd  132: out = 12'h408;
            14'd  133: out = 12'h408;
            14'd  134: out = 12'h408;
            14'd  135: out = 12'h409;
            14'd  136: out = 12'h409;
            14'd  137: out = 12'h409;
            14'd  138: out = 12'h409;
            14'd  139: out = 12'h409;
            14'd  140: out = 12'h409;
            14'd  141: out = 12'h409;
            14'd  142: out = 12'h409;
            14'd  143: out = 12'h409;
            14'd  144: out = 12'h409;
            14'd  145: out = 12'h409;
            14'd  146: out = 12'h409;
            14'd  147: out = 12'h409;
            14'd  148: out = 12'h409;
            14'd  149: out = 12'h409;
            14'd  150: out = 12'h409;
            14'd  151: out = 12'h40A;
            14'd  152: out = 12'h40A;
            14'd  153: out = 12'h40A;
            14'd  154: out = 12'h40A;
            14'd  155: out = 12'h40A;
            14'd  156: out = 12'h40A;
            14'd  157: out = 12'h40A;
            14'd  158: out = 12'h40A;
            14'd  159: out = 12'h40A;
            14'd  160: out = 12'h40A;
            14'd  161: out = 12'h40A;
            14'd  162: out = 12'h40A;
            14'd  163: out = 12'h40A;
            14'd  164: out = 12'h40A;
            14'd  165: out = 12'h40A;
            14'd  166: out = 12'h40A;
            14'd  167: out = 12'h40B;
            14'd  168: out = 12'h40B;
            14'd  169: out = 12'h40B;
            14'd  170: out = 12'h40B;
            14'd  171: out = 12'h40B;
            14'd  172: out = 12'h40B;
            14'd  173: out = 12'h40B;
            14'd  174: out = 12'h40B;
            14'd  175: out = 12'h40B;
            14'd  176: out = 12'h40B;
            14'd  177: out = 12'h40B;
            14'd  178: out = 12'h40B;
            14'd  179: out = 12'h40B;
            14'd  180: out = 12'h40B;
            14'd  181: out = 12'h40B;
            14'd  182: out = 12'h40C;
            14'd  183: out = 12'h40C;
            14'd  184: out = 12'h40C;
            14'd  185: out = 12'h40C;
            14'd  186: out = 12'h40C;
            14'd  187: out = 12'h40C;
            14'd  188: out = 12'h40C;
            14'd  189: out = 12'h40C;
            14'd  190: out = 12'h40C;
            14'd  191: out = 12'h40C;
            14'd  192: out = 12'h40C;
            14'd  193: out = 12'h40C;
            14'd  194: out = 12'h40C;
            14'd  195: out = 12'h40C;
            14'd  196: out = 12'h40C;
            14'd  197: out = 12'h40C;
            14'd  198: out = 12'h40D;
            14'd  199: out = 12'h40D;
            14'd  200: out = 12'h40D;
            14'd  201: out = 12'h40D;
            14'd  202: out = 12'h40D;
            14'd  203: out = 12'h40D;
            14'd  204: out = 12'h40D;
            14'd  205: out = 12'h40D;
            14'd  206: out = 12'h40D;
            14'd  207: out = 12'h40D;
            14'd  208: out = 12'h40D;
            14'd  209: out = 12'h40D;
            14'd  210: out = 12'h40D;
            14'd  211: out = 12'h40D;
            14'd  212: out = 12'h40D;
            14'd  213: out = 12'h40D;
            14'd  214: out = 12'h40E;
            14'd  215: out = 12'h40E;
            14'd  216: out = 12'h40E;
            14'd  217: out = 12'h40E;
            14'd  218: out = 12'h40E;
            14'd  219: out = 12'h40E;
            14'd  220: out = 12'h40E;
            14'd  221: out = 12'h40E;
            14'd  222: out = 12'h40E;
            14'd  223: out = 12'h40E;
            14'd  224: out = 12'h40E;
            14'd  225: out = 12'h40E;
            14'd  226: out = 12'h40E;
            14'd  227: out = 12'h40E;
            14'd  228: out = 12'h40E;
            14'd  229: out = 12'h40F;
            14'd  230: out = 12'h40F;
            14'd  231: out = 12'h40F;
            14'd  232: out = 12'h40F;
            14'd  233: out = 12'h40F;
            14'd  234: out = 12'h40F;
            14'd  235: out = 12'h40F;
            14'd  236: out = 12'h40F;
            14'd  237: out = 12'h40F;
            14'd  238: out = 12'h40F;
            14'd  239: out = 12'h40F;
            14'd  240: out = 12'h40F;
            14'd  241: out = 12'h40F;
            14'd  242: out = 12'h40F;
            14'd  243: out = 12'h40F;
            14'd  244: out = 12'h40F;
            14'd  245: out = 12'h410;
            14'd  246: out = 12'h410;
            14'd  247: out = 12'h410;
            14'd  248: out = 12'h410;
            14'd  249: out = 12'h410;
            14'd  250: out = 12'h410;
            14'd  251: out = 12'h410;
            14'd  252: out = 12'h410;
            14'd  253: out = 12'h410;
            14'd  254: out = 12'h410;
            14'd  255: out = 12'h410;
            14'd  256: out = 12'h410;
            14'd  257: out = 12'h410;
            14'd  258: out = 12'h410;
            14'd  259: out = 12'h410;
            14'd  260: out = 12'h411;
            14'd  261: out = 12'h411;
            14'd  262: out = 12'h411;
            14'd  263: out = 12'h411;
            14'd  264: out = 12'h411;
            14'd  265: out = 12'h411;
            14'd  266: out = 12'h411;
            14'd  267: out = 12'h411;
            14'd  268: out = 12'h411;
            14'd  269: out = 12'h411;
            14'd  270: out = 12'h411;
            14'd  271: out = 12'h411;
            14'd  272: out = 12'h411;
            14'd  273: out = 12'h411;
            14'd  274: out = 12'h411;
            14'd  275: out = 12'h411;
            14'd  276: out = 12'h412;
            14'd  277: out = 12'h412;
            14'd  278: out = 12'h412;
            14'd  279: out = 12'h412;
            14'd  280: out = 12'h412;
            14'd  281: out = 12'h412;
            14'd  282: out = 12'h412;
            14'd  283: out = 12'h412;
            14'd  284: out = 12'h412;
            14'd  285: out = 12'h412;
            14'd  286: out = 12'h412;
            14'd  287: out = 12'h412;
            14'd  288: out = 12'h412;
            14'd  289: out = 12'h412;
            14'd  290: out = 12'h412;
            14'd  291: out = 12'h413;
            14'd  292: out = 12'h413;
            14'd  293: out = 12'h413;
            14'd  294: out = 12'h413;
            14'd  295: out = 12'h413;
            14'd  296: out = 12'h413;
            14'd  297: out = 12'h413;
            14'd  298: out = 12'h413;
            14'd  299: out = 12'h413;
            14'd  300: out = 12'h413;
            14'd  301: out = 12'h413;
            14'd  302: out = 12'h413;
            14'd  303: out = 12'h413;
            14'd  304: out = 12'h413;
            14'd  305: out = 12'h413;
            14'd  306: out = 12'h413;
            14'd  307: out = 12'h414;
            14'd  308: out = 12'h414;
            14'd  309: out = 12'h414;
            14'd  310: out = 12'h414;
            14'd  311: out = 12'h414;
            14'd  312: out = 12'h414;
            14'd  313: out = 12'h414;
            14'd  314: out = 12'h414;
            14'd  315: out = 12'h414;
            14'd  316: out = 12'h414;
            14'd  317: out = 12'h414;
            14'd  318: out = 12'h414;
            14'd  319: out = 12'h414;
            14'd  320: out = 12'h414;
            14'd  321: out = 12'h414;
            14'd  322: out = 12'h415;
            14'd  323: out = 12'h415;
            14'd  324: out = 12'h415;
            14'd  325: out = 12'h415;
            14'd  326: out = 12'h415;
            14'd  327: out = 12'h415;
            14'd  328: out = 12'h415;
            14'd  329: out = 12'h415;
            14'd  330: out = 12'h415;
            14'd  331: out = 12'h415;
            14'd  332: out = 12'h415;
            14'd  333: out = 12'h415;
            14'd  334: out = 12'h415;
            14'd  335: out = 12'h415;
            14'd  336: out = 12'h415;
            14'd  337: out = 12'h416;
            14'd  338: out = 12'h416;
            14'd  339: out = 12'h416;
            14'd  340: out = 12'h416;
            14'd  341: out = 12'h416;
            14'd  342: out = 12'h416;
            14'd  343: out = 12'h416;
            14'd  344: out = 12'h416;
            14'd  345: out = 12'h416;
            14'd  346: out = 12'h416;
            14'd  347: out = 12'h416;
            14'd  348: out = 12'h416;
            14'd  349: out = 12'h416;
            14'd  350: out = 12'h416;
            14'd  351: out = 12'h416;
            14'd  352: out = 12'h416;
            14'd  353: out = 12'h417;
            14'd  354: out = 12'h417;
            14'd  355: out = 12'h417;
            14'd  356: out = 12'h417;
            14'd  357: out = 12'h417;
            14'd  358: out = 12'h417;
            14'd  359: out = 12'h417;
            14'd  360: out = 12'h417;
            14'd  361: out = 12'h417;
            14'd  362: out = 12'h417;
            14'd  363: out = 12'h417;
            14'd  364: out = 12'h417;
            14'd  365: out = 12'h417;
            14'd  366: out = 12'h417;
            14'd  367: out = 12'h417;
            14'd  368: out = 12'h418;
            14'd  369: out = 12'h418;
            14'd  370: out = 12'h418;
            14'd  371: out = 12'h418;
            14'd  372: out = 12'h418;
            14'd  373: out = 12'h418;
            14'd  374: out = 12'h418;
            14'd  375: out = 12'h418;
            14'd  376: out = 12'h418;
            14'd  377: out = 12'h418;
            14'd  378: out = 12'h418;
            14'd  379: out = 12'h418;
            14'd  380: out = 12'h418;
            14'd  381: out = 12'h418;
            14'd  382: out = 12'h418;
            14'd  383: out = 12'h419;
            14'd  384: out = 12'h419;
            14'd  385: out = 12'h419;
            14'd  386: out = 12'h419;
            14'd  387: out = 12'h419;
            14'd  388: out = 12'h419;
            14'd  389: out = 12'h419;
            14'd  390: out = 12'h419;
            14'd  391: out = 12'h419;
            14'd  392: out = 12'h419;
            14'd  393: out = 12'h419;
            14'd  394: out = 12'h419;
            14'd  395: out = 12'h419;
            14'd  396: out = 12'h419;
            14'd  397: out = 12'h419;
            14'd  398: out = 12'h419;
            14'd  399: out = 12'h41A;
            14'd  400: out = 12'h41A;
            14'd  401: out = 12'h41A;
            14'd  402: out = 12'h41A;
            14'd  403: out = 12'h41A;
            14'd  404: out = 12'h41A;
            14'd  405: out = 12'h41A;
            14'd  406: out = 12'h41A;
            14'd  407: out = 12'h41A;
            14'd  408: out = 12'h41A;
            14'd  409: out = 12'h41A;
            14'd  410: out = 12'h41A;
            14'd  411: out = 12'h41A;
            14'd  412: out = 12'h41A;
            14'd  413: out = 12'h41A;
            14'd  414: out = 12'h41B;
            14'd  415: out = 12'h41B;
            14'd  416: out = 12'h41B;
            14'd  417: out = 12'h41B;
            14'd  418: out = 12'h41B;
            14'd  419: out = 12'h41B;
            14'd  420: out = 12'h41B;
            14'd  421: out = 12'h41B;
            14'd  422: out = 12'h41B;
            14'd  423: out = 12'h41B;
            14'd  424: out = 12'h41B;
            14'd  425: out = 12'h41B;
            14'd  426: out = 12'h41B;
            14'd  427: out = 12'h41B;
            14'd  428: out = 12'h41B;
            14'd  429: out = 12'h41C;
            14'd  430: out = 12'h41C;
            14'd  431: out = 12'h41C;
            14'd  432: out = 12'h41C;
            14'd  433: out = 12'h41C;
            14'd  434: out = 12'h41C;
            14'd  435: out = 12'h41C;
            14'd  436: out = 12'h41C;
            14'd  437: out = 12'h41C;
            14'd  438: out = 12'h41C;
            14'd  439: out = 12'h41C;
            14'd  440: out = 12'h41C;
            14'd  441: out = 12'h41C;
            14'd  442: out = 12'h41C;
            14'd  443: out = 12'h41C;
            14'd  444: out = 12'h41D;
            14'd  445: out = 12'h41D;
            14'd  446: out = 12'h41D;
            14'd  447: out = 12'h41D;
            14'd  448: out = 12'h41D;
            14'd  449: out = 12'h41D;
            14'd  450: out = 12'h41D;
            14'd  451: out = 12'h41D;
            14'd  452: out = 12'h41D;
            14'd  453: out = 12'h41D;
            14'd  454: out = 12'h41D;
            14'd  455: out = 12'h41D;
            14'd  456: out = 12'h41D;
            14'd  457: out = 12'h41D;
            14'd  458: out = 12'h41D;
            14'd  459: out = 12'h41E;
            14'd  460: out = 12'h41E;
            14'd  461: out = 12'h41E;
            14'd  462: out = 12'h41E;
            14'd  463: out = 12'h41E;
            14'd  464: out = 12'h41E;
            14'd  465: out = 12'h41E;
            14'd  466: out = 12'h41E;
            14'd  467: out = 12'h41E;
            14'd  468: out = 12'h41E;
            14'd  469: out = 12'h41E;
            14'd  470: out = 12'h41E;
            14'd  471: out = 12'h41E;
            14'd  472: out = 12'h41E;
            14'd  473: out = 12'h41E;
            14'd  474: out = 12'h41F;
            14'd  475: out = 12'h41F;
            14'd  476: out = 12'h41F;
            14'd  477: out = 12'h41F;
            14'd  478: out = 12'h41F;
            14'd  479: out = 12'h41F;
            14'd  480: out = 12'h41F;
            14'd  481: out = 12'h41F;
            14'd  482: out = 12'h41F;
            14'd  483: out = 12'h41F;
            14'd  484: out = 12'h41F;
            14'd  485: out = 12'h41F;
            14'd  486: out = 12'h41F;
            14'd  487: out = 12'h41F;
            14'd  488: out = 12'h41F;
            14'd  489: out = 12'h420;
            14'd  490: out = 12'h420;
            14'd  491: out = 12'h420;
            14'd  492: out = 12'h420;
            14'd  493: out = 12'h420;
            14'd  494: out = 12'h420;
            14'd  495: out = 12'h420;
            14'd  496: out = 12'h420;
            14'd  497: out = 12'h420;
            14'd  498: out = 12'h420;
            14'd  499: out = 12'h420;
            14'd  500: out = 12'h420;
            14'd  501: out = 12'h420;
            14'd  502: out = 12'h420;
            14'd  503: out = 12'h420;
            14'd  504: out = 12'h420;
            14'd  505: out = 12'h421;
            14'd  506: out = 12'h421;
            14'd  507: out = 12'h421;
            14'd  508: out = 12'h421;
            14'd  509: out = 12'h421;
            14'd  510: out = 12'h421;
            14'd  511: out = 12'h421;
            14'd  512: out = 12'h421;
            14'd  513: out = 12'h421;
            14'd  514: out = 12'h421;
            14'd  515: out = 12'h421;
            14'd  516: out = 12'h421;
            14'd  517: out = 12'h421;
            14'd  518: out = 12'h421;
            14'd  519: out = 12'h421;
            14'd  520: out = 12'h422;
            14'd  521: out = 12'h422;
            14'd  522: out = 12'h422;
            14'd  523: out = 12'h422;
            14'd  524: out = 12'h422;
            14'd  525: out = 12'h422;
            14'd  526: out = 12'h422;
            14'd  527: out = 12'h422;
            14'd  528: out = 12'h422;
            14'd  529: out = 12'h422;
            14'd  530: out = 12'h422;
            14'd  531: out = 12'h422;
            14'd  532: out = 12'h422;
            14'd  533: out = 12'h422;
            14'd  534: out = 12'h422;
            14'd  535: out = 12'h423;
            14'd  536: out = 12'h423;
            14'd  537: out = 12'h423;
            14'd  538: out = 12'h423;
            14'd  539: out = 12'h423;
            14'd  540: out = 12'h423;
            14'd  541: out = 12'h423;
            14'd  542: out = 12'h423;
            14'd  543: out = 12'h423;
            14'd  544: out = 12'h423;
            14'd  545: out = 12'h423;
            14'd  546: out = 12'h423;
            14'd  547: out = 12'h423;
            14'd  548: out = 12'h423;
            14'd  549: out = 12'h424;
            14'd  550: out = 12'h424;
            14'd  551: out = 12'h424;
            14'd  552: out = 12'h424;
            14'd  553: out = 12'h424;
            14'd  554: out = 12'h424;
            14'd  555: out = 12'h424;
            14'd  556: out = 12'h424;
            14'd  557: out = 12'h424;
            14'd  558: out = 12'h424;
            14'd  559: out = 12'h424;
            14'd  560: out = 12'h424;
            14'd  561: out = 12'h424;
            14'd  562: out = 12'h424;
            14'd  563: out = 12'h424;
            14'd  564: out = 12'h425;
            14'd  565: out = 12'h425;
            14'd  566: out = 12'h425;
            14'd  567: out = 12'h425;
            14'd  568: out = 12'h425;
            14'd  569: out = 12'h425;
            14'd  570: out = 12'h425;
            14'd  571: out = 12'h425;
            14'd  572: out = 12'h425;
            14'd  573: out = 12'h425;
            14'd  574: out = 12'h425;
            14'd  575: out = 12'h425;
            14'd  576: out = 12'h425;
            14'd  577: out = 12'h425;
            14'd  578: out = 12'h425;
            14'd  579: out = 12'h426;
            14'd  580: out = 12'h426;
            14'd  581: out = 12'h426;
            14'd  582: out = 12'h426;
            14'd  583: out = 12'h426;
            14'd  584: out = 12'h426;
            14'd  585: out = 12'h426;
            14'd  586: out = 12'h426;
            14'd  587: out = 12'h426;
            14'd  588: out = 12'h426;
            14'd  589: out = 12'h426;
            14'd  590: out = 12'h426;
            14'd  591: out = 12'h426;
            14'd  592: out = 12'h426;
            14'd  593: out = 12'h426;
            14'd  594: out = 12'h427;
            14'd  595: out = 12'h427;
            14'd  596: out = 12'h427;
            14'd  597: out = 12'h427;
            14'd  598: out = 12'h427;
            14'd  599: out = 12'h427;
            14'd  600: out = 12'h427;
            14'd  601: out = 12'h427;
            14'd  602: out = 12'h427;
            14'd  603: out = 12'h427;
            14'd  604: out = 12'h427;
            14'd  605: out = 12'h427;
            14'd  606: out = 12'h427;
            14'd  607: out = 12'h427;
            14'd  608: out = 12'h427;
            14'd  609: out = 12'h428;
            14'd  610: out = 12'h428;
            14'd  611: out = 12'h428;
            14'd  612: out = 12'h428;
            14'd  613: out = 12'h428;
            14'd  614: out = 12'h428;
            14'd  615: out = 12'h428;
            14'd  616: out = 12'h428;
            14'd  617: out = 12'h428;
            14'd  618: out = 12'h428;
            14'd  619: out = 12'h428;
            14'd  620: out = 12'h428;
            14'd  621: out = 12'h428;
            14'd  622: out = 12'h428;
            14'd  623: out = 12'h428;
            14'd  624: out = 12'h429;
            14'd  625: out = 12'h429;
            14'd  626: out = 12'h429;
            14'd  627: out = 12'h429;
            14'd  628: out = 12'h429;
            14'd  629: out = 12'h429;
            14'd  630: out = 12'h429;
            14'd  631: out = 12'h429;
            14'd  632: out = 12'h429;
            14'd  633: out = 12'h429;
            14'd  634: out = 12'h429;
            14'd  635: out = 12'h429;
            14'd  636: out = 12'h429;
            14'd  637: out = 12'h429;
            14'd  638: out = 12'h429;
            14'd  639: out = 12'h42A;
            14'd  640: out = 12'h42A;
            14'd  641: out = 12'h42A;
            14'd  642: out = 12'h42A;
            14'd  643: out = 12'h42A;
            14'd  644: out = 12'h42A;
            14'd  645: out = 12'h42A;
            14'd  646: out = 12'h42A;
            14'd  647: out = 12'h42A;
            14'd  648: out = 12'h42A;
            14'd  649: out = 12'h42A;
            14'd  650: out = 12'h42A;
            14'd  651: out = 12'h42A;
            14'd  652: out = 12'h42A;
            14'd  653: out = 12'h42B;
            14'd  654: out = 12'h42B;
            14'd  655: out = 12'h42B;
            14'd  656: out = 12'h42B;
            14'd  657: out = 12'h42B;
            14'd  658: out = 12'h42B;
            14'd  659: out = 12'h42B;
            14'd  660: out = 12'h42B;
            14'd  661: out = 12'h42B;
            14'd  662: out = 12'h42B;
            14'd  663: out = 12'h42B;
            14'd  664: out = 12'h42B;
            14'd  665: out = 12'h42B;
            14'd  666: out = 12'h42B;
            14'd  667: out = 12'h42B;
            14'd  668: out = 12'h42C;
            14'd  669: out = 12'h42C;
            14'd  670: out = 12'h42C;
            14'd  671: out = 12'h42C;
            14'd  672: out = 12'h42C;
            14'd  673: out = 12'h42C;
            14'd  674: out = 12'h42C;
            14'd  675: out = 12'h42C;
            14'd  676: out = 12'h42C;
            14'd  677: out = 12'h42C;
            14'd  678: out = 12'h42C;
            14'd  679: out = 12'h42C;
            14'd  680: out = 12'h42C;
            14'd  681: out = 12'h42C;
            14'd  682: out = 12'h42C;
            14'd  683: out = 12'h42D;
            14'd  684: out = 12'h42D;
            14'd  685: out = 12'h42D;
            14'd  686: out = 12'h42D;
            14'd  687: out = 12'h42D;
            14'd  688: out = 12'h42D;
            14'd  689: out = 12'h42D;
            14'd  690: out = 12'h42D;
            14'd  691: out = 12'h42D;
            14'd  692: out = 12'h42D;
            14'd  693: out = 12'h42D;
            14'd  694: out = 12'h42D;
            14'd  695: out = 12'h42D;
            14'd  696: out = 12'h42D;
            14'd  697: out = 12'h42D;
            14'd  698: out = 12'h42E;
            14'd  699: out = 12'h42E;
            14'd  700: out = 12'h42E;
            14'd  701: out = 12'h42E;
            14'd  702: out = 12'h42E;
            14'd  703: out = 12'h42E;
            14'd  704: out = 12'h42E;
            14'd  705: out = 12'h42E;
            14'd  706: out = 12'h42E;
            14'd  707: out = 12'h42E;
            14'd  708: out = 12'h42E;
            14'd  709: out = 12'h42E;
            14'd  710: out = 12'h42E;
            14'd  711: out = 12'h42E;
            14'd  712: out = 12'h42F;
            14'd  713: out = 12'h42F;
            14'd  714: out = 12'h42F;
            14'd  715: out = 12'h42F;
            14'd  716: out = 12'h42F;
            14'd  717: out = 12'h42F;
            14'd  718: out = 12'h42F;
            14'd  719: out = 12'h42F;
            14'd  720: out = 12'h42F;
            14'd  721: out = 12'h42F;
            14'd  722: out = 12'h42F;
            14'd  723: out = 12'h42F;
            14'd  724: out = 12'h42F;
            14'd  725: out = 12'h42F;
            14'd  726: out = 12'h42F;
            14'd  727: out = 12'h430;
            14'd  728: out = 12'h430;
            14'd  729: out = 12'h430;
            14'd  730: out = 12'h430;
            14'd  731: out = 12'h430;
            14'd  732: out = 12'h430;
            14'd  733: out = 12'h430;
            14'd  734: out = 12'h430;
            14'd  735: out = 12'h430;
            14'd  736: out = 12'h430;
            14'd  737: out = 12'h430;
            14'd  738: out = 12'h430;
            14'd  739: out = 12'h430;
            14'd  740: out = 12'h430;
            14'd  741: out = 12'h431;
            14'd  742: out = 12'h431;
            14'd  743: out = 12'h431;
            14'd  744: out = 12'h431;
            14'd  745: out = 12'h431;
            14'd  746: out = 12'h431;
            14'd  747: out = 12'h431;
            14'd  748: out = 12'h431;
            14'd  749: out = 12'h431;
            14'd  750: out = 12'h431;
            14'd  751: out = 12'h431;
            14'd  752: out = 12'h431;
            14'd  753: out = 12'h431;
            14'd  754: out = 12'h431;
            14'd  755: out = 12'h431;
            14'd  756: out = 12'h432;
            14'd  757: out = 12'h432;
            14'd  758: out = 12'h432;
            14'd  759: out = 12'h432;
            14'd  760: out = 12'h432;
            14'd  761: out = 12'h432;
            14'd  762: out = 12'h432;
            14'd  763: out = 12'h432;
            14'd  764: out = 12'h432;
            14'd  765: out = 12'h432;
            14'd  766: out = 12'h432;
            14'd  767: out = 12'h432;
            14'd  768: out = 12'h432;
            14'd  769: out = 12'h432;
            14'd  770: out = 12'h432;
            14'd  771: out = 12'h433;
            14'd  772: out = 12'h433;
            14'd  773: out = 12'h433;
            14'd  774: out = 12'h433;
            14'd  775: out = 12'h433;
            14'd  776: out = 12'h433;
            14'd  777: out = 12'h433;
            14'd  778: out = 12'h433;
            14'd  779: out = 12'h433;
            14'd  780: out = 12'h433;
            14'd  781: out = 12'h433;
            14'd  782: out = 12'h433;
            14'd  783: out = 12'h433;
            14'd  784: out = 12'h433;
            14'd  785: out = 12'h434;
            14'd  786: out = 12'h434;
            14'd  787: out = 12'h434;
            14'd  788: out = 12'h434;
            14'd  789: out = 12'h434;
            14'd  790: out = 12'h434;
            14'd  791: out = 12'h434;
            14'd  792: out = 12'h434;
            14'd  793: out = 12'h434;
            14'd  794: out = 12'h434;
            14'd  795: out = 12'h434;
            14'd  796: out = 12'h434;
            14'd  797: out = 12'h434;
            14'd  798: out = 12'h434;
            14'd  799: out = 12'h434;
            14'd  800: out = 12'h435;
            14'd  801: out = 12'h435;
            14'd  802: out = 12'h435;
            14'd  803: out = 12'h435;
            14'd  804: out = 12'h435;
            14'd  805: out = 12'h435;
            14'd  806: out = 12'h435;
            14'd  807: out = 12'h435;
            14'd  808: out = 12'h435;
            14'd  809: out = 12'h435;
            14'd  810: out = 12'h435;
            14'd  811: out = 12'h435;
            14'd  812: out = 12'h435;
            14'd  813: out = 12'h435;
            14'd  814: out = 12'h436;
            14'd  815: out = 12'h436;
            14'd  816: out = 12'h436;
            14'd  817: out = 12'h436;
            14'd  818: out = 12'h436;
            14'd  819: out = 12'h436;
            14'd  820: out = 12'h436;
            14'd  821: out = 12'h436;
            14'd  822: out = 12'h436;
            14'd  823: out = 12'h436;
            14'd  824: out = 12'h436;
            14'd  825: out = 12'h436;
            14'd  826: out = 12'h436;
            14'd  827: out = 12'h436;
            14'd  828: out = 12'h437;
            14'd  829: out = 12'h437;
            14'd  830: out = 12'h437;
            14'd  831: out = 12'h437;
            14'd  832: out = 12'h437;
            14'd  833: out = 12'h437;
            14'd  834: out = 12'h437;
            14'd  835: out = 12'h437;
            14'd  836: out = 12'h437;
            14'd  837: out = 12'h437;
            14'd  838: out = 12'h437;
            14'd  839: out = 12'h437;
            14'd  840: out = 12'h437;
            14'd  841: out = 12'h437;
            14'd  842: out = 12'h437;
            14'd  843: out = 12'h438;
            14'd  844: out = 12'h438;
            14'd  845: out = 12'h438;
            14'd  846: out = 12'h438;
            14'd  847: out = 12'h438;
            14'd  848: out = 12'h438;
            14'd  849: out = 12'h438;
            14'd  850: out = 12'h438;
            14'd  851: out = 12'h438;
            14'd  852: out = 12'h438;
            14'd  853: out = 12'h438;
            14'd  854: out = 12'h438;
            14'd  855: out = 12'h438;
            14'd  856: out = 12'h438;
            14'd  857: out = 12'h439;
            14'd  858: out = 12'h439;
            14'd  859: out = 12'h439;
            14'd  860: out = 12'h439;
            14'd  861: out = 12'h439;
            14'd  862: out = 12'h439;
            14'd  863: out = 12'h439;
            14'd  864: out = 12'h439;
            14'd  865: out = 12'h439;
            14'd  866: out = 12'h439;
            14'd  867: out = 12'h439;
            14'd  868: out = 12'h439;
            14'd  869: out = 12'h439;
            14'd  870: out = 12'h439;
            14'd  871: out = 12'h439;
            14'd  872: out = 12'h43A;
            14'd  873: out = 12'h43A;
            14'd  874: out = 12'h43A;
            14'd  875: out = 12'h43A;
            14'd  876: out = 12'h43A;
            14'd  877: out = 12'h43A;
            14'd  878: out = 12'h43A;
            14'd  879: out = 12'h43A;
            14'd  880: out = 12'h43A;
            14'd  881: out = 12'h43A;
            14'd  882: out = 12'h43A;
            14'd  883: out = 12'h43A;
            14'd  884: out = 12'h43A;
            14'd  885: out = 12'h43A;
            14'd  886: out = 12'h43B;
            14'd  887: out = 12'h43B;
            14'd  888: out = 12'h43B;
            14'd  889: out = 12'h43B;
            14'd  890: out = 12'h43B;
            14'd  891: out = 12'h43B;
            14'd  892: out = 12'h43B;
            14'd  893: out = 12'h43B;
            14'd  894: out = 12'h43B;
            14'd  895: out = 12'h43B;
            14'd  896: out = 12'h43B;
            14'd  897: out = 12'h43B;
            14'd  898: out = 12'h43B;
            14'd  899: out = 12'h43B;
            14'd  900: out = 12'h43C;
            14'd  901: out = 12'h43C;
            14'd  902: out = 12'h43C;
            14'd  903: out = 12'h43C;
            14'd  904: out = 12'h43C;
            14'd  905: out = 12'h43C;
            14'd  906: out = 12'h43C;
            14'd  907: out = 12'h43C;
            14'd  908: out = 12'h43C;
            14'd  909: out = 12'h43C;
            14'd  910: out = 12'h43C;
            14'd  911: out = 12'h43C;
            14'd  912: out = 12'h43C;
            14'd  913: out = 12'h43C;
            14'd  914: out = 12'h43D;
            14'd  915: out = 12'h43D;
            14'd  916: out = 12'h43D;
            14'd  917: out = 12'h43D;
            14'd  918: out = 12'h43D;
            14'd  919: out = 12'h43D;
            14'd  920: out = 12'h43D;
            14'd  921: out = 12'h43D;
            14'd  922: out = 12'h43D;
            14'd  923: out = 12'h43D;
            14'd  924: out = 12'h43D;
            14'd  925: out = 12'h43D;
            14'd  926: out = 12'h43D;
            14'd  927: out = 12'h43D;
            14'd  928: out = 12'h43D;
            14'd  929: out = 12'h43E;
            14'd  930: out = 12'h43E;
            14'd  931: out = 12'h43E;
            14'd  932: out = 12'h43E;
            14'd  933: out = 12'h43E;
            14'd  934: out = 12'h43E;
            14'd  935: out = 12'h43E;
            14'd  936: out = 12'h43E;
            14'd  937: out = 12'h43E;
            14'd  938: out = 12'h43E;
            14'd  939: out = 12'h43E;
            14'd  940: out = 12'h43E;
            14'd  941: out = 12'h43E;
            14'd  942: out = 12'h43E;
            14'd  943: out = 12'h43F;
            14'd  944: out = 12'h43F;
            14'd  945: out = 12'h43F;
            14'd  946: out = 12'h43F;
            14'd  947: out = 12'h43F;
            14'd  948: out = 12'h43F;
            14'd  949: out = 12'h43F;
            14'd  950: out = 12'h43F;
            14'd  951: out = 12'h43F;
            14'd  952: out = 12'h43F;
            14'd  953: out = 12'h43F;
            14'd  954: out = 12'h43F;
            14'd  955: out = 12'h43F;
            14'd  956: out = 12'h43F;
            14'd  957: out = 12'h440;
            14'd  958: out = 12'h440;
            14'd  959: out = 12'h440;
            14'd  960: out = 12'h440;
            14'd  961: out = 12'h440;
            14'd  962: out = 12'h440;
            14'd  963: out = 12'h440;
            14'd  964: out = 12'h440;
            14'd  965: out = 12'h440;
            14'd  966: out = 12'h440;
            14'd  967: out = 12'h440;
            14'd  968: out = 12'h440;
            14'd  969: out = 12'h440;
            14'd  970: out = 12'h440;
            14'd  971: out = 12'h441;
            14'd  972: out = 12'h441;
            14'd  973: out = 12'h441;
            14'd  974: out = 12'h441;
            14'd  975: out = 12'h441;
            14'd  976: out = 12'h441;
            14'd  977: out = 12'h441;
            14'd  978: out = 12'h441;
            14'd  979: out = 12'h441;
            14'd  980: out = 12'h441;
            14'd  981: out = 12'h441;
            14'd  982: out = 12'h441;
            14'd  983: out = 12'h441;
            14'd  984: out = 12'h441;
            14'd  985: out = 12'h442;
            14'd  986: out = 12'h442;
            14'd  987: out = 12'h442;
            14'd  988: out = 12'h442;
            14'd  989: out = 12'h442;
            14'd  990: out = 12'h442;
            14'd  991: out = 12'h442;
            14'd  992: out = 12'h442;
            14'd  993: out = 12'h442;
            14'd  994: out = 12'h442;
            14'd  995: out = 12'h442;
            14'd  996: out = 12'h442;
            14'd  997: out = 12'h442;
            14'd  998: out = 12'h442;
            14'd  999: out = 12'h442;
            14'd 1000: out = 12'h443;
            14'd 1001: out = 12'h443;
            14'd 1002: out = 12'h443;
            14'd 1003: out = 12'h443;
            14'd 1004: out = 12'h443;
            14'd 1005: out = 12'h443;
            14'd 1006: out = 12'h443;
            14'd 1007: out = 12'h443;
            14'd 1008: out = 12'h443;
            14'd 1009: out = 12'h443;
            14'd 1010: out = 12'h443;
            14'd 1011: out = 12'h443;
            14'd 1012: out = 12'h443;
            14'd 1013: out = 12'h443;
            14'd 1014: out = 12'h444;
            14'd 1015: out = 12'h444;
            14'd 1016: out = 12'h444;
            14'd 1017: out = 12'h444;
            14'd 1018: out = 12'h444;
            14'd 1019: out = 12'h444;
            14'd 1020: out = 12'h444;
            14'd 1021: out = 12'h444;
            14'd 1022: out = 12'h444;
            14'd 1023: out = 12'h444;
            14'd 1024: out = 12'h444;
            14'd 1025: out = 12'h444;
            14'd 1026: out = 12'h444;
            14'd 1027: out = 12'h444;
            14'd 1028: out = 12'h445;
            14'd 1029: out = 12'h445;
            14'd 1030: out = 12'h445;
            14'd 1031: out = 12'h445;
            14'd 1032: out = 12'h445;
            14'd 1033: out = 12'h445;
            14'd 1034: out = 12'h445;
            14'd 1035: out = 12'h445;
            14'd 1036: out = 12'h445;
            14'd 1037: out = 12'h445;
            14'd 1038: out = 12'h445;
            14'd 1039: out = 12'h445;
            14'd 1040: out = 12'h445;
            14'd 1041: out = 12'h445;
            14'd 1042: out = 12'h446;
            14'd 1043: out = 12'h446;
            14'd 1044: out = 12'h446;
            14'd 1045: out = 12'h446;
            14'd 1046: out = 12'h446;
            14'd 1047: out = 12'h446;
            14'd 1048: out = 12'h446;
            14'd 1049: out = 12'h446;
            14'd 1050: out = 12'h446;
            14'd 1051: out = 12'h446;
            14'd 1052: out = 12'h446;
            14'd 1053: out = 12'h446;
            14'd 1054: out = 12'h446;
            14'd 1055: out = 12'h446;
            14'd 1056: out = 12'h447;
            14'd 1057: out = 12'h447;
            14'd 1058: out = 12'h447;
            14'd 1059: out = 12'h447;
            14'd 1060: out = 12'h447;
            14'd 1061: out = 12'h447;
            14'd 1062: out = 12'h447;
            14'd 1063: out = 12'h447;
            14'd 1064: out = 12'h447;
            14'd 1065: out = 12'h447;
            14'd 1066: out = 12'h447;
            14'd 1067: out = 12'h447;
            14'd 1068: out = 12'h447;
            14'd 1069: out = 12'h447;
            14'd 1070: out = 12'h448;
            14'd 1071: out = 12'h448;
            14'd 1072: out = 12'h448;
            14'd 1073: out = 12'h448;
            14'd 1074: out = 12'h448;
            14'd 1075: out = 12'h448;
            14'd 1076: out = 12'h448;
            14'd 1077: out = 12'h448;
            14'd 1078: out = 12'h448;
            14'd 1079: out = 12'h448;
            14'd 1080: out = 12'h448;
            14'd 1081: out = 12'h448;
            14'd 1082: out = 12'h448;
            14'd 1083: out = 12'h448;
            14'd 1084: out = 12'h449;
            14'd 1085: out = 12'h449;
            14'd 1086: out = 12'h449;
            14'd 1087: out = 12'h449;
            14'd 1088: out = 12'h449;
            14'd 1089: out = 12'h449;
            14'd 1090: out = 12'h449;
            14'd 1091: out = 12'h449;
            14'd 1092: out = 12'h449;
            14'd 1093: out = 12'h449;
            14'd 1094: out = 12'h449;
            14'd 1095: out = 12'h449;
            14'd 1096: out = 12'h449;
            14'd 1097: out = 12'h449;
            14'd 1098: out = 12'h44A;
            14'd 1099: out = 12'h44A;
            14'd 1100: out = 12'h44A;
            14'd 1101: out = 12'h44A;
            14'd 1102: out = 12'h44A;
            14'd 1103: out = 12'h44A;
            14'd 1104: out = 12'h44A;
            14'd 1105: out = 12'h44A;
            14'd 1106: out = 12'h44A;
            14'd 1107: out = 12'h44A;
            14'd 1108: out = 12'h44A;
            14'd 1109: out = 12'h44A;
            14'd 1110: out = 12'h44A;
            14'd 1111: out = 12'h44A;
            14'd 1112: out = 12'h44B;
            14'd 1113: out = 12'h44B;
            14'd 1114: out = 12'h44B;
            14'd 1115: out = 12'h44B;
            14'd 1116: out = 12'h44B;
            14'd 1117: out = 12'h44B;
            14'd 1118: out = 12'h44B;
            14'd 1119: out = 12'h44B;
            14'd 1120: out = 12'h44B;
            14'd 1121: out = 12'h44B;
            14'd 1122: out = 12'h44B;
            14'd 1123: out = 12'h44B;
            14'd 1124: out = 12'h44B;
            14'd 1125: out = 12'h44B;
            14'd 1126: out = 12'h44C;
            14'd 1127: out = 12'h44C;
            14'd 1128: out = 12'h44C;
            14'd 1129: out = 12'h44C;
            14'd 1130: out = 12'h44C;
            14'd 1131: out = 12'h44C;
            14'd 1132: out = 12'h44C;
            14'd 1133: out = 12'h44C;
            14'd 1134: out = 12'h44C;
            14'd 1135: out = 12'h44C;
            14'd 1136: out = 12'h44C;
            14'd 1137: out = 12'h44C;
            14'd 1138: out = 12'h44C;
            14'd 1139: out = 12'h44D;
            14'd 1140: out = 12'h44D;
            14'd 1141: out = 12'h44D;
            14'd 1142: out = 12'h44D;
            14'd 1143: out = 12'h44D;
            14'd 1144: out = 12'h44D;
            14'd 1145: out = 12'h44D;
            14'd 1146: out = 12'h44D;
            14'd 1147: out = 12'h44D;
            14'd 1148: out = 12'h44D;
            14'd 1149: out = 12'h44D;
            14'd 1150: out = 12'h44D;
            14'd 1151: out = 12'h44D;
            14'd 1152: out = 12'h44D;
            14'd 1153: out = 12'h44E;
            14'd 1154: out = 12'h44E;
            14'd 1155: out = 12'h44E;
            14'd 1156: out = 12'h44E;
            14'd 1157: out = 12'h44E;
            14'd 1158: out = 12'h44E;
            14'd 1159: out = 12'h44E;
            14'd 1160: out = 12'h44E;
            14'd 1161: out = 12'h44E;
            14'd 1162: out = 12'h44E;
            14'd 1163: out = 12'h44E;
            14'd 1164: out = 12'h44E;
            14'd 1165: out = 12'h44E;
            14'd 1166: out = 12'h44E;
            14'd 1167: out = 12'h44F;
            14'd 1168: out = 12'h44F;
            14'd 1169: out = 12'h44F;
            14'd 1170: out = 12'h44F;
            14'd 1171: out = 12'h44F;
            14'd 1172: out = 12'h44F;
            14'd 1173: out = 12'h44F;
            14'd 1174: out = 12'h44F;
            14'd 1175: out = 12'h44F;
            14'd 1176: out = 12'h44F;
            14'd 1177: out = 12'h44F;
            14'd 1178: out = 12'h44F;
            14'd 1179: out = 12'h44F;
            14'd 1180: out = 12'h44F;
            14'd 1181: out = 12'h450;
            14'd 1182: out = 12'h450;
            14'd 1183: out = 12'h450;
            14'd 1184: out = 12'h450;
            14'd 1185: out = 12'h450;
            14'd 1186: out = 12'h450;
            14'd 1187: out = 12'h450;
            14'd 1188: out = 12'h450;
            14'd 1189: out = 12'h450;
            14'd 1190: out = 12'h450;
            14'd 1191: out = 12'h450;
            14'd 1192: out = 12'h450;
            14'd 1193: out = 12'h450;
            14'd 1194: out = 12'h450;
            14'd 1195: out = 12'h451;
            14'd 1196: out = 12'h451;
            14'd 1197: out = 12'h451;
            14'd 1198: out = 12'h451;
            14'd 1199: out = 12'h451;
            14'd 1200: out = 12'h451;
            14'd 1201: out = 12'h451;
            14'd 1202: out = 12'h451;
            14'd 1203: out = 12'h451;
            14'd 1204: out = 12'h451;
            14'd 1205: out = 12'h451;
            14'd 1206: out = 12'h451;
            14'd 1207: out = 12'h451;
            14'd 1208: out = 12'h452;
            14'd 1209: out = 12'h452;
            14'd 1210: out = 12'h452;
            14'd 1211: out = 12'h452;
            14'd 1212: out = 12'h452;
            14'd 1213: out = 12'h452;
            14'd 1214: out = 12'h452;
            14'd 1215: out = 12'h452;
            14'd 1216: out = 12'h452;
            14'd 1217: out = 12'h452;
            14'd 1218: out = 12'h452;
            14'd 1219: out = 12'h452;
            14'd 1220: out = 12'h452;
            14'd 1221: out = 12'h452;
            14'd 1222: out = 12'h453;
            14'd 1223: out = 12'h453;
            14'd 1224: out = 12'h453;
            14'd 1225: out = 12'h453;
            14'd 1226: out = 12'h453;
            14'd 1227: out = 12'h453;
            14'd 1228: out = 12'h453;
            14'd 1229: out = 12'h453;
            14'd 1230: out = 12'h453;
            14'd 1231: out = 12'h453;
            14'd 1232: out = 12'h453;
            14'd 1233: out = 12'h453;
            14'd 1234: out = 12'h453;
            14'd 1235: out = 12'h453;
            14'd 1236: out = 12'h454;
            14'd 1237: out = 12'h454;
            14'd 1238: out = 12'h454;
            14'd 1239: out = 12'h454;
            14'd 1240: out = 12'h454;
            14'd 1241: out = 12'h454;
            14'd 1242: out = 12'h454;
            14'd 1243: out = 12'h454;
            14'd 1244: out = 12'h454;
            14'd 1245: out = 12'h454;
            14'd 1246: out = 12'h454;
            14'd 1247: out = 12'h454;
            14'd 1248: out = 12'h454;
            14'd 1249: out = 12'h455;
            14'd 1250: out = 12'h455;
            14'd 1251: out = 12'h455;
            14'd 1252: out = 12'h455;
            14'd 1253: out = 12'h455;
            14'd 1254: out = 12'h455;
            14'd 1255: out = 12'h455;
            14'd 1256: out = 12'h455;
            14'd 1257: out = 12'h455;
            14'd 1258: out = 12'h455;
            14'd 1259: out = 12'h455;
            14'd 1260: out = 12'h455;
            14'd 1261: out = 12'h455;
            14'd 1262: out = 12'h455;
            14'd 1263: out = 12'h456;
            14'd 1264: out = 12'h456;
            14'd 1265: out = 12'h456;
            14'd 1266: out = 12'h456;
            14'd 1267: out = 12'h456;
            14'd 1268: out = 12'h456;
            14'd 1269: out = 12'h456;
            14'd 1270: out = 12'h456;
            14'd 1271: out = 12'h456;
            14'd 1272: out = 12'h456;
            14'd 1273: out = 12'h456;
            14'd 1274: out = 12'h456;
            14'd 1275: out = 12'h456;
            14'd 1276: out = 12'h456;
            14'd 1277: out = 12'h457;
            14'd 1278: out = 12'h457;
            14'd 1279: out = 12'h457;
            14'd 1280: out = 12'h457;
            14'd 1281: out = 12'h457;
            14'd 1282: out = 12'h457;
            14'd 1283: out = 12'h457;
            14'd 1284: out = 12'h457;
            14'd 1285: out = 12'h457;
            14'd 1286: out = 12'h457;
            14'd 1287: out = 12'h457;
            14'd 1288: out = 12'h457;
            14'd 1289: out = 12'h457;
            14'd 1290: out = 12'h458;
            14'd 1291: out = 12'h458;
            14'd 1292: out = 12'h458;
            14'd 1293: out = 12'h458;
            14'd 1294: out = 12'h458;
            14'd 1295: out = 12'h458;
            14'd 1296: out = 12'h458;
            14'd 1297: out = 12'h458;
            14'd 1298: out = 12'h458;
            14'd 1299: out = 12'h458;
            14'd 1300: out = 12'h458;
            14'd 1301: out = 12'h458;
            14'd 1302: out = 12'h458;
            14'd 1303: out = 12'h458;
            14'd 1304: out = 12'h459;
            14'd 1305: out = 12'h459;
            14'd 1306: out = 12'h459;
            14'd 1307: out = 12'h459;
            14'd 1308: out = 12'h459;
            14'd 1309: out = 12'h459;
            14'd 1310: out = 12'h459;
            14'd 1311: out = 12'h459;
            14'd 1312: out = 12'h459;
            14'd 1313: out = 12'h459;
            14'd 1314: out = 12'h459;
            14'd 1315: out = 12'h459;
            14'd 1316: out = 12'h459;
            14'd 1317: out = 12'h45A;
            14'd 1318: out = 12'h45A;
            14'd 1319: out = 12'h45A;
            14'd 1320: out = 12'h45A;
            14'd 1321: out = 12'h45A;
            14'd 1322: out = 12'h45A;
            14'd 1323: out = 12'h45A;
            14'd 1324: out = 12'h45A;
            14'd 1325: out = 12'h45A;
            14'd 1326: out = 12'h45A;
            14'd 1327: out = 12'h45A;
            14'd 1328: out = 12'h45A;
            14'd 1329: out = 12'h45A;
            14'd 1330: out = 12'h45A;
            14'd 1331: out = 12'h45B;
            14'd 1332: out = 12'h45B;
            14'd 1333: out = 12'h45B;
            14'd 1334: out = 12'h45B;
            14'd 1335: out = 12'h45B;
            14'd 1336: out = 12'h45B;
            14'd 1337: out = 12'h45B;
            14'd 1338: out = 12'h45B;
            14'd 1339: out = 12'h45B;
            14'd 1340: out = 12'h45B;
            14'd 1341: out = 12'h45B;
            14'd 1342: out = 12'h45B;
            14'd 1343: out = 12'h45B;
            14'd 1344: out = 12'h45C;
            14'd 1345: out = 12'h45C;
            14'd 1346: out = 12'h45C;
            14'd 1347: out = 12'h45C;
            14'd 1348: out = 12'h45C;
            14'd 1349: out = 12'h45C;
            14'd 1350: out = 12'h45C;
            14'd 1351: out = 12'h45C;
            14'd 1352: out = 12'h45C;
            14'd 1353: out = 12'h45C;
            14'd 1354: out = 12'h45C;
            14'd 1355: out = 12'h45C;
            14'd 1356: out = 12'h45C;
            14'd 1357: out = 12'h45C;
            14'd 1358: out = 12'h45D;
            14'd 1359: out = 12'h45D;
            14'd 1360: out = 12'h45D;
            14'd 1361: out = 12'h45D;
            14'd 1362: out = 12'h45D;
            14'd 1363: out = 12'h45D;
            14'd 1364: out = 12'h45D;
            14'd 1365: out = 12'h45D;
            14'd 1366: out = 12'h45D;
            14'd 1367: out = 12'h45D;
            14'd 1368: out = 12'h45D;
            14'd 1369: out = 12'h45D;
            14'd 1370: out = 12'h45D;
            14'd 1371: out = 12'h45E;
            14'd 1372: out = 12'h45E;
            14'd 1373: out = 12'h45E;
            14'd 1374: out = 12'h45E;
            14'd 1375: out = 12'h45E;
            14'd 1376: out = 12'h45E;
            14'd 1377: out = 12'h45E;
            14'd 1378: out = 12'h45E;
            14'd 1379: out = 12'h45E;
            14'd 1380: out = 12'h45E;
            14'd 1381: out = 12'h45E;
            14'd 1382: out = 12'h45E;
            14'd 1383: out = 12'h45E;
            14'd 1384: out = 12'h45E;
            14'd 1385: out = 12'h45F;
            14'd 1386: out = 12'h45F;
            14'd 1387: out = 12'h45F;
            14'd 1388: out = 12'h45F;
            14'd 1389: out = 12'h45F;
            14'd 1390: out = 12'h45F;
            14'd 1391: out = 12'h45F;
            14'd 1392: out = 12'h45F;
            14'd 1393: out = 12'h45F;
            14'd 1394: out = 12'h45F;
            14'd 1395: out = 12'h45F;
            14'd 1396: out = 12'h45F;
            14'd 1397: out = 12'h45F;
            14'd 1398: out = 12'h460;
            14'd 1399: out = 12'h460;
            14'd 1400: out = 12'h460;
            14'd 1401: out = 12'h460;
            14'd 1402: out = 12'h460;
            14'd 1403: out = 12'h460;
            14'd 1404: out = 12'h460;
            14'd 1405: out = 12'h460;
            14'd 1406: out = 12'h460;
            14'd 1407: out = 12'h460;
            14'd 1408: out = 12'h460;
            14'd 1409: out = 12'h460;
            14'd 1410: out = 12'h460;
            14'd 1411: out = 12'h460;
            14'd 1412: out = 12'h461;
            14'd 1413: out = 12'h461;
            14'd 1414: out = 12'h461;
            14'd 1415: out = 12'h461;
            14'd 1416: out = 12'h461;
            14'd 1417: out = 12'h461;
            14'd 1418: out = 12'h461;
            14'd 1419: out = 12'h461;
            14'd 1420: out = 12'h461;
            14'd 1421: out = 12'h461;
            14'd 1422: out = 12'h461;
            14'd 1423: out = 12'h461;
            14'd 1424: out = 12'h461;
            14'd 1425: out = 12'h462;
            14'd 1426: out = 12'h462;
            14'd 1427: out = 12'h462;
            14'd 1428: out = 12'h462;
            14'd 1429: out = 12'h462;
            14'd 1430: out = 12'h462;
            14'd 1431: out = 12'h462;
            14'd 1432: out = 12'h462;
            14'd 1433: out = 12'h462;
            14'd 1434: out = 12'h462;
            14'd 1435: out = 12'h462;
            14'd 1436: out = 12'h462;
            14'd 1437: out = 12'h462;
            14'd 1438: out = 12'h463;
            14'd 1439: out = 12'h463;
            14'd 1440: out = 12'h463;
            14'd 1441: out = 12'h463;
            14'd 1442: out = 12'h463;
            14'd 1443: out = 12'h463;
            14'd 1444: out = 12'h463;
            14'd 1445: out = 12'h463;
            14'd 1446: out = 12'h463;
            14'd 1447: out = 12'h463;
            14'd 1448: out = 12'h463;
            14'd 1449: out = 12'h463;
            14'd 1450: out = 12'h463;
            14'd 1451: out = 12'h463;
            14'd 1452: out = 12'h464;
            14'd 1453: out = 12'h464;
            14'd 1454: out = 12'h464;
            14'd 1455: out = 12'h464;
            14'd 1456: out = 12'h464;
            14'd 1457: out = 12'h464;
            14'd 1458: out = 12'h464;
            14'd 1459: out = 12'h464;
            14'd 1460: out = 12'h464;
            14'd 1461: out = 12'h464;
            14'd 1462: out = 12'h464;
            14'd 1463: out = 12'h464;
            14'd 1464: out = 12'h464;
            14'd 1465: out = 12'h465;
            14'd 1466: out = 12'h465;
            14'd 1467: out = 12'h465;
            14'd 1468: out = 12'h465;
            14'd 1469: out = 12'h465;
            14'd 1470: out = 12'h465;
            14'd 1471: out = 12'h465;
            14'd 1472: out = 12'h465;
            14'd 1473: out = 12'h465;
            14'd 1474: out = 12'h465;
            14'd 1475: out = 12'h465;
            14'd 1476: out = 12'h465;
            14'd 1477: out = 12'h465;
            14'd 1478: out = 12'h466;
            14'd 1479: out = 12'h466;
            14'd 1480: out = 12'h466;
            14'd 1481: out = 12'h466;
            14'd 1482: out = 12'h466;
            14'd 1483: out = 12'h466;
            14'd 1484: out = 12'h466;
            14'd 1485: out = 12'h466;
            14'd 1486: out = 12'h466;
            14'd 1487: out = 12'h466;
            14'd 1488: out = 12'h466;
            14'd 1489: out = 12'h466;
            14'd 1490: out = 12'h466;
            14'd 1491: out = 12'h467;
            14'd 1492: out = 12'h467;
            14'd 1493: out = 12'h467;
            14'd 1494: out = 12'h467;
            14'd 1495: out = 12'h467;
            14'd 1496: out = 12'h467;
            14'd 1497: out = 12'h467;
            14'd 1498: out = 12'h467;
            14'd 1499: out = 12'h467;
            14'd 1500: out = 12'h467;
            14'd 1501: out = 12'h467;
            14'd 1502: out = 12'h467;
            14'd 1503: out = 12'h467;
            14'd 1504: out = 12'h468;
            14'd 1505: out = 12'h468;
            14'd 1506: out = 12'h468;
            14'd 1507: out = 12'h468;
            14'd 1508: out = 12'h468;
            14'd 1509: out = 12'h468;
            14'd 1510: out = 12'h468;
            14'd 1511: out = 12'h468;
            14'd 1512: out = 12'h468;
            14'd 1513: out = 12'h468;
            14'd 1514: out = 12'h468;
            14'd 1515: out = 12'h468;
            14'd 1516: out = 12'h468;
            14'd 1517: out = 12'h468;
            14'd 1518: out = 12'h469;
            14'd 1519: out = 12'h469;
            14'd 1520: out = 12'h469;
            14'd 1521: out = 12'h469;
            14'd 1522: out = 12'h469;
            14'd 1523: out = 12'h469;
            14'd 1524: out = 12'h469;
            14'd 1525: out = 12'h469;
            14'd 1526: out = 12'h469;
            14'd 1527: out = 12'h469;
            14'd 1528: out = 12'h469;
            14'd 1529: out = 12'h469;
            14'd 1530: out = 12'h469;
            14'd 1531: out = 12'h46A;
            14'd 1532: out = 12'h46A;
            14'd 1533: out = 12'h46A;
            14'd 1534: out = 12'h46A;
            14'd 1535: out = 12'h46A;
            14'd 1536: out = 12'h46A;
            14'd 1537: out = 12'h46A;
            14'd 1538: out = 12'h46A;
            14'd 1539: out = 12'h46A;
            14'd 1540: out = 12'h46A;
            14'd 1541: out = 12'h46A;
            14'd 1542: out = 12'h46A;
            14'd 1543: out = 12'h46A;
            14'd 1544: out = 12'h46B;
            14'd 1545: out = 12'h46B;
            14'd 1546: out = 12'h46B;
            14'd 1547: out = 12'h46B;
            14'd 1548: out = 12'h46B;
            14'd 1549: out = 12'h46B;
            14'd 1550: out = 12'h46B;
            14'd 1551: out = 12'h46B;
            14'd 1552: out = 12'h46B;
            14'd 1553: out = 12'h46B;
            14'd 1554: out = 12'h46B;
            14'd 1555: out = 12'h46B;
            14'd 1556: out = 12'h46B;
            14'd 1557: out = 12'h46C;
            14'd 1558: out = 12'h46C;
            14'd 1559: out = 12'h46C;
            14'd 1560: out = 12'h46C;
            14'd 1561: out = 12'h46C;
            14'd 1562: out = 12'h46C;
            14'd 1563: out = 12'h46C;
            14'd 1564: out = 12'h46C;
            14'd 1565: out = 12'h46C;
            14'd 1566: out = 12'h46C;
            14'd 1567: out = 12'h46C;
            14'd 1568: out = 12'h46C;
            14'd 1569: out = 12'h46C;
            14'd 1570: out = 12'h46D;
            14'd 1571: out = 12'h46D;
            14'd 1572: out = 12'h46D;
            14'd 1573: out = 12'h46D;
            14'd 1574: out = 12'h46D;
            14'd 1575: out = 12'h46D;
            14'd 1576: out = 12'h46D;
            14'd 1577: out = 12'h46D;
            14'd 1578: out = 12'h46D;
            14'd 1579: out = 12'h46D;
            14'd 1580: out = 12'h46D;
            14'd 1581: out = 12'h46D;
            14'd 1582: out = 12'h46D;
            14'd 1583: out = 12'h46E;
            14'd 1584: out = 12'h46E;
            14'd 1585: out = 12'h46E;
            14'd 1586: out = 12'h46E;
            14'd 1587: out = 12'h46E;
            14'd 1588: out = 12'h46E;
            14'd 1589: out = 12'h46E;
            14'd 1590: out = 12'h46E;
            14'd 1591: out = 12'h46E;
            14'd 1592: out = 12'h46E;
            14'd 1593: out = 12'h46E;
            14'd 1594: out = 12'h46E;
            14'd 1595: out = 12'h46E;
            14'd 1596: out = 12'h46F;
            14'd 1597: out = 12'h46F;
            14'd 1598: out = 12'h46F;
            14'd 1599: out = 12'h46F;
            14'd 1600: out = 12'h46F;
            14'd 1601: out = 12'h46F;
            14'd 1602: out = 12'h46F;
            14'd 1603: out = 12'h46F;
            14'd 1604: out = 12'h46F;
            14'd 1605: out = 12'h46F;
            14'd 1606: out = 12'h46F;
            14'd 1607: out = 12'h46F;
            14'd 1608: out = 12'h46F;
            14'd 1609: out = 12'h470;
            14'd 1610: out = 12'h470;
            14'd 1611: out = 12'h470;
            14'd 1612: out = 12'h470;
            14'd 1613: out = 12'h470;
            14'd 1614: out = 12'h470;
            14'd 1615: out = 12'h470;
            14'd 1616: out = 12'h470;
            14'd 1617: out = 12'h470;
            14'd 1618: out = 12'h470;
            14'd 1619: out = 12'h470;
            14'd 1620: out = 12'h470;
            14'd 1621: out = 12'h470;
            14'd 1622: out = 12'h471;
            14'd 1623: out = 12'h471;
            14'd 1624: out = 12'h471;
            14'd 1625: out = 12'h471;
            14'd 1626: out = 12'h471;
            14'd 1627: out = 12'h471;
            14'd 1628: out = 12'h471;
            14'd 1629: out = 12'h471;
            14'd 1630: out = 12'h471;
            14'd 1631: out = 12'h471;
            14'd 1632: out = 12'h471;
            14'd 1633: out = 12'h471;
            14'd 1634: out = 12'h471;
            14'd 1635: out = 12'h472;
            14'd 1636: out = 12'h472;
            14'd 1637: out = 12'h472;
            14'd 1638: out = 12'h472;
            14'd 1639: out = 12'h472;
            14'd 1640: out = 12'h472;
            14'd 1641: out = 12'h472;
            14'd 1642: out = 12'h472;
            14'd 1643: out = 12'h472;
            14'd 1644: out = 12'h472;
            14'd 1645: out = 12'h472;
            14'd 1646: out = 12'h472;
            14'd 1647: out = 12'h472;
            14'd 1648: out = 12'h473;
            14'd 1649: out = 12'h473;
            14'd 1650: out = 12'h473;
            14'd 1651: out = 12'h473;
            14'd 1652: out = 12'h473;
            14'd 1653: out = 12'h473;
            14'd 1654: out = 12'h473;
            14'd 1655: out = 12'h473;
            14'd 1656: out = 12'h473;
            14'd 1657: out = 12'h473;
            14'd 1658: out = 12'h473;
            14'd 1659: out = 12'h473;
            14'd 1660: out = 12'h473;
            14'd 1661: out = 12'h474;
            14'd 1662: out = 12'h474;
            14'd 1663: out = 12'h474;
            14'd 1664: out = 12'h474;
            14'd 1665: out = 12'h474;
            14'd 1666: out = 12'h474;
            14'd 1667: out = 12'h474;
            14'd 1668: out = 12'h474;
            14'd 1669: out = 12'h474;
            14'd 1670: out = 12'h474;
            14'd 1671: out = 12'h474;
            14'd 1672: out = 12'h474;
            14'd 1673: out = 12'h474;
            14'd 1674: out = 12'h475;
            14'd 1675: out = 12'h475;
            14'd 1676: out = 12'h475;
            14'd 1677: out = 12'h475;
            14'd 1678: out = 12'h475;
            14'd 1679: out = 12'h475;
            14'd 1680: out = 12'h475;
            14'd 1681: out = 12'h475;
            14'd 1682: out = 12'h475;
            14'd 1683: out = 12'h475;
            14'd 1684: out = 12'h475;
            14'd 1685: out = 12'h475;
            14'd 1686: out = 12'h475;
            14'd 1687: out = 12'h476;
            14'd 1688: out = 12'h476;
            14'd 1689: out = 12'h476;
            14'd 1690: out = 12'h476;
            14'd 1691: out = 12'h476;
            14'd 1692: out = 12'h476;
            14'd 1693: out = 12'h476;
            14'd 1694: out = 12'h476;
            14'd 1695: out = 12'h476;
            14'd 1696: out = 12'h476;
            14'd 1697: out = 12'h476;
            14'd 1698: out = 12'h476;
            14'd 1699: out = 12'h476;
            14'd 1700: out = 12'h477;
            14'd 1701: out = 12'h477;
            14'd 1702: out = 12'h477;
            14'd 1703: out = 12'h477;
            14'd 1704: out = 12'h477;
            14'd 1705: out = 12'h477;
            14'd 1706: out = 12'h477;
            14'd 1707: out = 12'h477;
            14'd 1708: out = 12'h477;
            14'd 1709: out = 12'h477;
            14'd 1710: out = 12'h477;
            14'd 1711: out = 12'h477;
            14'd 1712: out = 12'h477;
            14'd 1713: out = 12'h478;
            14'd 1714: out = 12'h478;
            14'd 1715: out = 12'h478;
            14'd 1716: out = 12'h478;
            14'd 1717: out = 12'h478;
            14'd 1718: out = 12'h478;
            14'd 1719: out = 12'h478;
            14'd 1720: out = 12'h478;
            14'd 1721: out = 12'h478;
            14'd 1722: out = 12'h478;
            14'd 1723: out = 12'h478;
            14'd 1724: out = 12'h478;
            14'd 1725: out = 12'h478;
            14'd 1726: out = 12'h479;
            14'd 1727: out = 12'h479;
            14'd 1728: out = 12'h479;
            14'd 1729: out = 12'h479;
            14'd 1730: out = 12'h479;
            14'd 1731: out = 12'h479;
            14'd 1732: out = 12'h479;
            14'd 1733: out = 12'h479;
            14'd 1734: out = 12'h479;
            14'd 1735: out = 12'h479;
            14'd 1736: out = 12'h479;
            14'd 1737: out = 12'h479;
            14'd 1738: out = 12'h47A;
            14'd 1739: out = 12'h47A;
            14'd 1740: out = 12'h47A;
            14'd 1741: out = 12'h47A;
            14'd 1742: out = 12'h47A;
            14'd 1743: out = 12'h47A;
            14'd 1744: out = 12'h47A;
            14'd 1745: out = 12'h47A;
            14'd 1746: out = 12'h47A;
            14'd 1747: out = 12'h47A;
            14'd 1748: out = 12'h47A;
            14'd 1749: out = 12'h47A;
            14'd 1750: out = 12'h47A;
            14'd 1751: out = 12'h47B;
            14'd 1752: out = 12'h47B;
            14'd 1753: out = 12'h47B;
            14'd 1754: out = 12'h47B;
            14'd 1755: out = 12'h47B;
            14'd 1756: out = 12'h47B;
            14'd 1757: out = 12'h47B;
            14'd 1758: out = 12'h47B;
            14'd 1759: out = 12'h47B;
            14'd 1760: out = 12'h47B;
            14'd 1761: out = 12'h47B;
            14'd 1762: out = 12'h47B;
            14'd 1763: out = 12'h47B;
            14'd 1764: out = 12'h47C;
            14'd 1765: out = 12'h47C;
            14'd 1766: out = 12'h47C;
            14'd 1767: out = 12'h47C;
            14'd 1768: out = 12'h47C;
            14'd 1769: out = 12'h47C;
            14'd 1770: out = 12'h47C;
            14'd 1771: out = 12'h47C;
            14'd 1772: out = 12'h47C;
            14'd 1773: out = 12'h47C;
            14'd 1774: out = 12'h47C;
            14'd 1775: out = 12'h47C;
            14'd 1776: out = 12'h47C;
            14'd 1777: out = 12'h47D;
            14'd 1778: out = 12'h47D;
            14'd 1779: out = 12'h47D;
            14'd 1780: out = 12'h47D;
            14'd 1781: out = 12'h47D;
            14'd 1782: out = 12'h47D;
            14'd 1783: out = 12'h47D;
            14'd 1784: out = 12'h47D;
            14'd 1785: out = 12'h47D;
            14'd 1786: out = 12'h47D;
            14'd 1787: out = 12'h47D;
            14'd 1788: out = 12'h47D;
            14'd 1789: out = 12'h47E;
            14'd 1790: out = 12'h47E;
            14'd 1791: out = 12'h47E;
            14'd 1792: out = 12'h47E;
            14'd 1793: out = 12'h47E;
            14'd 1794: out = 12'h47E;
            14'd 1795: out = 12'h47E;
            14'd 1796: out = 12'h47E;
            14'd 1797: out = 12'h47E;
            14'd 1798: out = 12'h47E;
            14'd 1799: out = 12'h47E;
            14'd 1800: out = 12'h47E;
            14'd 1801: out = 12'h47E;
            14'd 1802: out = 12'h47F;
            14'd 1803: out = 12'h47F;
            14'd 1804: out = 12'h47F;
            14'd 1805: out = 12'h47F;
            14'd 1806: out = 12'h47F;
            14'd 1807: out = 12'h47F;
            14'd 1808: out = 12'h47F;
            14'd 1809: out = 12'h47F;
            14'd 1810: out = 12'h47F;
            14'd 1811: out = 12'h47F;
            14'd 1812: out = 12'h47F;
            14'd 1813: out = 12'h47F;
            14'd 1814: out = 12'h47F;
            14'd 1815: out = 12'h480;
            14'd 1816: out = 12'h480;
            14'd 1817: out = 12'h480;
            14'd 1818: out = 12'h480;
            14'd 1819: out = 12'h480;
            14'd 1820: out = 12'h480;
            14'd 1821: out = 12'h480;
            14'd 1822: out = 12'h480;
            14'd 1823: out = 12'h480;
            14'd 1824: out = 12'h480;
            14'd 1825: out = 12'h480;
            14'd 1826: out = 12'h480;
            14'd 1827: out = 12'h481;
            14'd 1828: out = 12'h481;
            14'd 1829: out = 12'h481;
            14'd 1830: out = 12'h481;
            14'd 1831: out = 12'h481;
            14'd 1832: out = 12'h481;
            14'd 1833: out = 12'h481;
            14'd 1834: out = 12'h481;
            14'd 1835: out = 12'h481;
            14'd 1836: out = 12'h481;
            14'd 1837: out = 12'h481;
            14'd 1838: out = 12'h481;
            14'd 1839: out = 12'h481;
            14'd 1840: out = 12'h482;
            14'd 1841: out = 12'h482;
            14'd 1842: out = 12'h482;
            14'd 1843: out = 12'h482;
            14'd 1844: out = 12'h482;
            14'd 1845: out = 12'h482;
            14'd 1846: out = 12'h482;
            14'd 1847: out = 12'h482;
            14'd 1848: out = 12'h482;
            14'd 1849: out = 12'h482;
            14'd 1850: out = 12'h482;
            14'd 1851: out = 12'h482;
            14'd 1852: out = 12'h483;
            14'd 1853: out = 12'h483;
            14'd 1854: out = 12'h483;
            14'd 1855: out = 12'h483;
            14'd 1856: out = 12'h483;
            14'd 1857: out = 12'h483;
            14'd 1858: out = 12'h483;
            14'd 1859: out = 12'h483;
            14'd 1860: out = 12'h483;
            14'd 1861: out = 12'h483;
            14'd 1862: out = 12'h483;
            14'd 1863: out = 12'h483;
            14'd 1864: out = 12'h483;
            14'd 1865: out = 12'h484;
            14'd 1866: out = 12'h484;
            14'd 1867: out = 12'h484;
            14'd 1868: out = 12'h484;
            14'd 1869: out = 12'h484;
            14'd 1870: out = 12'h484;
            14'd 1871: out = 12'h484;
            14'd 1872: out = 12'h484;
            14'd 1873: out = 12'h484;
            14'd 1874: out = 12'h484;
            14'd 1875: out = 12'h484;
            14'd 1876: out = 12'h484;
            14'd 1877: out = 12'h484;
            14'd 1878: out = 12'h485;
            14'd 1879: out = 12'h485;
            14'd 1880: out = 12'h485;
            14'd 1881: out = 12'h485;
            14'd 1882: out = 12'h485;
            14'd 1883: out = 12'h485;
            14'd 1884: out = 12'h485;
            14'd 1885: out = 12'h485;
            14'd 1886: out = 12'h485;
            14'd 1887: out = 12'h485;
            14'd 1888: out = 12'h485;
            14'd 1889: out = 12'h485;
            14'd 1890: out = 12'h486;
            14'd 1891: out = 12'h486;
            14'd 1892: out = 12'h486;
            14'd 1893: out = 12'h486;
            14'd 1894: out = 12'h486;
            14'd 1895: out = 12'h486;
            14'd 1896: out = 12'h486;
            14'd 1897: out = 12'h486;
            14'd 1898: out = 12'h486;
            14'd 1899: out = 12'h486;
            14'd 1900: out = 12'h486;
            14'd 1901: out = 12'h486;
            14'd 1902: out = 12'h486;
            14'd 1903: out = 12'h487;
            14'd 1904: out = 12'h487;
            14'd 1905: out = 12'h487;
            14'd 1906: out = 12'h487;
            14'd 1907: out = 12'h487;
            14'd 1908: out = 12'h487;
            14'd 1909: out = 12'h487;
            14'd 1910: out = 12'h487;
            14'd 1911: out = 12'h487;
            14'd 1912: out = 12'h487;
            14'd 1913: out = 12'h487;
            14'd 1914: out = 12'h487;
            14'd 1915: out = 12'h488;
            14'd 1916: out = 12'h488;
            14'd 1917: out = 12'h488;
            14'd 1918: out = 12'h488;
            14'd 1919: out = 12'h488;
            14'd 1920: out = 12'h488;
            14'd 1921: out = 12'h488;
            14'd 1922: out = 12'h488;
            14'd 1923: out = 12'h488;
            14'd 1924: out = 12'h488;
            14'd 1925: out = 12'h488;
            14'd 1926: out = 12'h488;
            14'd 1927: out = 12'h488;
            14'd 1928: out = 12'h489;
            14'd 1929: out = 12'h489;
            14'd 1930: out = 12'h489;
            14'd 1931: out = 12'h489;
            14'd 1932: out = 12'h489;
            14'd 1933: out = 12'h489;
            14'd 1934: out = 12'h489;
            14'd 1935: out = 12'h489;
            14'd 1936: out = 12'h489;
            14'd 1937: out = 12'h489;
            14'd 1938: out = 12'h489;
            14'd 1939: out = 12'h489;
            14'd 1940: out = 12'h48A;
            14'd 1941: out = 12'h48A;
            14'd 1942: out = 12'h48A;
            14'd 1943: out = 12'h48A;
            14'd 1944: out = 12'h48A;
            14'd 1945: out = 12'h48A;
            14'd 1946: out = 12'h48A;
            14'd 1947: out = 12'h48A;
            14'd 1948: out = 12'h48A;
            14'd 1949: out = 12'h48A;
            14'd 1950: out = 12'h48A;
            14'd 1951: out = 12'h48A;
            14'd 1952: out = 12'h48B;
            14'd 1953: out = 12'h48B;
            14'd 1954: out = 12'h48B;
            14'd 1955: out = 12'h48B;
            14'd 1956: out = 12'h48B;
            14'd 1957: out = 12'h48B;
            14'd 1958: out = 12'h48B;
            14'd 1959: out = 12'h48B;
            14'd 1960: out = 12'h48B;
            14'd 1961: out = 12'h48B;
            14'd 1962: out = 12'h48B;
            14'd 1963: out = 12'h48B;
            14'd 1964: out = 12'h48B;
            14'd 1965: out = 12'h48C;
            14'd 1966: out = 12'h48C;
            14'd 1967: out = 12'h48C;
            14'd 1968: out = 12'h48C;
            14'd 1969: out = 12'h48C;
            14'd 1970: out = 12'h48C;
            14'd 1971: out = 12'h48C;
            14'd 1972: out = 12'h48C;
            14'd 1973: out = 12'h48C;
            14'd 1974: out = 12'h48C;
            14'd 1975: out = 12'h48C;
            14'd 1976: out = 12'h48C;
            14'd 1977: out = 12'h48D;
            14'd 1978: out = 12'h48D;
            14'd 1979: out = 12'h48D;
            14'd 1980: out = 12'h48D;
            14'd 1981: out = 12'h48D;
            14'd 1982: out = 12'h48D;
            14'd 1983: out = 12'h48D;
            14'd 1984: out = 12'h48D;
            14'd 1985: out = 12'h48D;
            14'd 1986: out = 12'h48D;
            14'd 1987: out = 12'h48D;
            14'd 1988: out = 12'h48D;
            14'd 1989: out = 12'h48D;
            14'd 1990: out = 12'h48E;
            14'd 1991: out = 12'h48E;
            14'd 1992: out = 12'h48E;
            14'd 1993: out = 12'h48E;
            14'd 1994: out = 12'h48E;
            14'd 1995: out = 12'h48E;
            14'd 1996: out = 12'h48E;
            14'd 1997: out = 12'h48E;
            14'd 1998: out = 12'h48E;
            14'd 1999: out = 12'h48E;
            14'd 2000: out = 12'h48E;
            14'd 2001: out = 12'h48E;
            14'd 2002: out = 12'h48F;
            14'd 2003: out = 12'h48F;
            14'd 2004: out = 12'h48F;
            14'd 2005: out = 12'h48F;
            14'd 2006: out = 12'h48F;
            14'd 2007: out = 12'h48F;
            14'd 2008: out = 12'h48F;
            14'd 2009: out = 12'h48F;
            14'd 2010: out = 12'h48F;
            14'd 2011: out = 12'h48F;
            14'd 2012: out = 12'h48F;
            14'd 2013: out = 12'h48F;
            14'd 2014: out = 12'h490;
            14'd 2015: out = 12'h490;
            14'd 2016: out = 12'h490;
            14'd 2017: out = 12'h490;
            14'd 2018: out = 12'h490;
            14'd 2019: out = 12'h490;
            14'd 2020: out = 12'h490;
            14'd 2021: out = 12'h490;
            14'd 2022: out = 12'h490;
            14'd 2023: out = 12'h490;
            14'd 2024: out = 12'h490;
            14'd 2025: out = 12'h490;
            14'd 2026: out = 12'h490;
            14'd 2027: out = 12'h491;
            14'd 2028: out = 12'h491;
            14'd 2029: out = 12'h491;
            14'd 2030: out = 12'h491;
            14'd 2031: out = 12'h491;
            14'd 2032: out = 12'h491;
            14'd 2033: out = 12'h491;
            14'd 2034: out = 12'h491;
            14'd 2035: out = 12'h491;
            14'd 2036: out = 12'h491;
            14'd 2037: out = 12'h491;
            14'd 2038: out = 12'h491;
            14'd 2039: out = 12'h492;
            14'd 2040: out = 12'h492;
            14'd 2041: out = 12'h492;
            14'd 2042: out = 12'h492;
            14'd 2043: out = 12'h492;
            14'd 2044: out = 12'h492;
            14'd 2045: out = 12'h492;
            14'd 2046: out = 12'h492;
            14'd 2047: out = 12'h492;
            14'd 2048: out = 12'h492;
            14'd 2049: out = 12'h492;
            14'd 2050: out = 12'h492;
            14'd 2051: out = 12'h493;
            14'd 2052: out = 12'h493;
            14'd 2053: out = 12'h493;
            14'd 2054: out = 12'h493;
            14'd 2055: out = 12'h493;
            14'd 2056: out = 12'h493;
            14'd 2057: out = 12'h493;
            14'd 2058: out = 12'h493;
            14'd 2059: out = 12'h493;
            14'd 2060: out = 12'h493;
            14'd 2061: out = 12'h493;
            14'd 2062: out = 12'h493;
            14'd 2063: out = 12'h494;
            14'd 2064: out = 12'h494;
            14'd 2065: out = 12'h494;
            14'd 2066: out = 12'h494;
            14'd 2067: out = 12'h494;
            14'd 2068: out = 12'h494;
            14'd 2069: out = 12'h494;
            14'd 2070: out = 12'h494;
            14'd 2071: out = 12'h494;
            14'd 2072: out = 12'h494;
            14'd 2073: out = 12'h494;
            14'd 2074: out = 12'h494;
            14'd 2075: out = 12'h494;
            14'd 2076: out = 12'h495;
            14'd 2077: out = 12'h495;
            14'd 2078: out = 12'h495;
            14'd 2079: out = 12'h495;
            14'd 2080: out = 12'h495;
            14'd 2081: out = 12'h495;
            14'd 2082: out = 12'h495;
            14'd 2083: out = 12'h495;
            14'd 2084: out = 12'h495;
            14'd 2085: out = 12'h495;
            14'd 2086: out = 12'h495;
            14'd 2087: out = 12'h495;
            14'd 2088: out = 12'h496;
            14'd 2089: out = 12'h496;
            14'd 2090: out = 12'h496;
            14'd 2091: out = 12'h496;
            14'd 2092: out = 12'h496;
            14'd 2093: out = 12'h496;
            14'd 2094: out = 12'h496;
            14'd 2095: out = 12'h496;
            14'd 2096: out = 12'h496;
            14'd 2097: out = 12'h496;
            14'd 2098: out = 12'h496;
            14'd 2099: out = 12'h496;
            14'd 2100: out = 12'h497;
            14'd 2101: out = 12'h497;
            14'd 2102: out = 12'h497;
            14'd 2103: out = 12'h497;
            14'd 2104: out = 12'h497;
            14'd 2105: out = 12'h497;
            14'd 2106: out = 12'h497;
            14'd 2107: out = 12'h497;
            14'd 2108: out = 12'h497;
            14'd 2109: out = 12'h497;
            14'd 2110: out = 12'h497;
            14'd 2111: out = 12'h497;
            14'd 2112: out = 12'h498;
            14'd 2113: out = 12'h498;
            14'd 2114: out = 12'h498;
            14'd 2115: out = 12'h498;
            14'd 2116: out = 12'h498;
            14'd 2117: out = 12'h498;
            14'd 2118: out = 12'h498;
            14'd 2119: out = 12'h498;
            14'd 2120: out = 12'h498;
            14'd 2121: out = 12'h498;
            14'd 2122: out = 12'h498;
            14'd 2123: out = 12'h498;
            14'd 2124: out = 12'h499;
            14'd 2125: out = 12'h499;
            14'd 2126: out = 12'h499;
            14'd 2127: out = 12'h499;
            14'd 2128: out = 12'h499;
            14'd 2129: out = 12'h499;
            14'd 2130: out = 12'h499;
            14'd 2131: out = 12'h499;
            14'd 2132: out = 12'h499;
            14'd 2133: out = 12'h499;
            14'd 2134: out = 12'h499;
            14'd 2135: out = 12'h499;
            14'd 2136: out = 12'h49A;
            14'd 2137: out = 12'h49A;
            14'd 2138: out = 12'h49A;
            14'd 2139: out = 12'h49A;
            14'd 2140: out = 12'h49A;
            14'd 2141: out = 12'h49A;
            14'd 2142: out = 12'h49A;
            14'd 2143: out = 12'h49A;
            14'd 2144: out = 12'h49A;
            14'd 2145: out = 12'h49A;
            14'd 2146: out = 12'h49A;
            14'd 2147: out = 12'h49A;
            14'd 2148: out = 12'h49B;
            14'd 2149: out = 12'h49B;
            14'd 2150: out = 12'h49B;
            14'd 2151: out = 12'h49B;
            14'd 2152: out = 12'h49B;
            14'd 2153: out = 12'h49B;
            14'd 2154: out = 12'h49B;
            14'd 2155: out = 12'h49B;
            14'd 2156: out = 12'h49B;
            14'd 2157: out = 12'h49B;
            14'd 2158: out = 12'h49B;
            14'd 2159: out = 12'h49B;
            14'd 2160: out = 12'h49C;
            14'd 2161: out = 12'h49C;
            14'd 2162: out = 12'h49C;
            14'd 2163: out = 12'h49C;
            14'd 2164: out = 12'h49C;
            14'd 2165: out = 12'h49C;
            14'd 2166: out = 12'h49C;
            14'd 2167: out = 12'h49C;
            14'd 2168: out = 12'h49C;
            14'd 2169: out = 12'h49C;
            14'd 2170: out = 12'h49C;
            14'd 2171: out = 12'h49C;
            14'd 2172: out = 12'h49C;
            14'd 2173: out = 12'h49D;
            14'd 2174: out = 12'h49D;
            14'd 2175: out = 12'h49D;
            14'd 2176: out = 12'h49D;
            14'd 2177: out = 12'h49D;
            14'd 2178: out = 12'h49D;
            14'd 2179: out = 12'h49D;
            14'd 2180: out = 12'h49D;
            14'd 2181: out = 12'h49D;
            14'd 2182: out = 12'h49D;
            14'd 2183: out = 12'h49D;
            14'd 2184: out = 12'h49D;
            14'd 2185: out = 12'h49E;
            14'd 2186: out = 12'h49E;
            14'd 2187: out = 12'h49E;
            14'd 2188: out = 12'h49E;
            14'd 2189: out = 12'h49E;
            14'd 2190: out = 12'h49E;
            14'd 2191: out = 12'h49E;
            14'd 2192: out = 12'h49E;
            14'd 2193: out = 12'h49E;
            14'd 2194: out = 12'h49E;
            14'd 2195: out = 12'h49E;
            14'd 2196: out = 12'h49E;
            14'd 2197: out = 12'h49F;
            14'd 2198: out = 12'h49F;
            14'd 2199: out = 12'h49F;
            14'd 2200: out = 12'h49F;
            14'd 2201: out = 12'h49F;
            14'd 2202: out = 12'h49F;
            14'd 2203: out = 12'h49F;
            14'd 2204: out = 12'h49F;
            14'd 2205: out = 12'h49F;
            14'd 2206: out = 12'h49F;
            14'd 2207: out = 12'h49F;
            14'd 2208: out = 12'h49F;
            14'd 2209: out = 12'h4A0;
            14'd 2210: out = 12'h4A0;
            14'd 2211: out = 12'h4A0;
            14'd 2212: out = 12'h4A0;
            14'd 2213: out = 12'h4A0;
            14'd 2214: out = 12'h4A0;
            14'd 2215: out = 12'h4A0;
            14'd 2216: out = 12'h4A0;
            14'd 2217: out = 12'h4A0;
            14'd 2218: out = 12'h4A0;
            14'd 2219: out = 12'h4A0;
            14'd 2220: out = 12'h4A0;
            14'd 2221: out = 12'h4A1;
            14'd 2222: out = 12'h4A1;
            14'd 2223: out = 12'h4A1;
            14'd 2224: out = 12'h4A1;
            14'd 2225: out = 12'h4A1;
            14'd 2226: out = 12'h4A1;
            14'd 2227: out = 12'h4A1;
            14'd 2228: out = 12'h4A1;
            14'd 2229: out = 12'h4A1;
            14'd 2230: out = 12'h4A1;
            14'd 2231: out = 12'h4A1;
            14'd 2232: out = 12'h4A2;
            14'd 2233: out = 12'h4A2;
            14'd 2234: out = 12'h4A2;
            14'd 2235: out = 12'h4A2;
            14'd 2236: out = 12'h4A2;
            14'd 2237: out = 12'h4A2;
            14'd 2238: out = 12'h4A2;
            14'd 2239: out = 12'h4A2;
            14'd 2240: out = 12'h4A2;
            14'd 2241: out = 12'h4A2;
            14'd 2242: out = 12'h4A2;
            14'd 2243: out = 12'h4A2;
            14'd 2244: out = 12'h4A3;
            14'd 2245: out = 12'h4A3;
            14'd 2246: out = 12'h4A3;
            14'd 2247: out = 12'h4A3;
            14'd 2248: out = 12'h4A3;
            14'd 2249: out = 12'h4A3;
            14'd 2250: out = 12'h4A3;
            14'd 2251: out = 12'h4A3;
            14'd 2252: out = 12'h4A3;
            14'd 2253: out = 12'h4A3;
            14'd 2254: out = 12'h4A3;
            14'd 2255: out = 12'h4A3;
            14'd 2256: out = 12'h4A4;
            14'd 2257: out = 12'h4A4;
            14'd 2258: out = 12'h4A4;
            14'd 2259: out = 12'h4A4;
            14'd 2260: out = 12'h4A4;
            14'd 2261: out = 12'h4A4;
            14'd 2262: out = 12'h4A4;
            14'd 2263: out = 12'h4A4;
            14'd 2264: out = 12'h4A4;
            14'd 2265: out = 12'h4A4;
            14'd 2266: out = 12'h4A4;
            14'd 2267: out = 12'h4A4;
            14'd 2268: out = 12'h4A5;
            14'd 2269: out = 12'h4A5;
            14'd 2270: out = 12'h4A5;
            14'd 2271: out = 12'h4A5;
            14'd 2272: out = 12'h4A5;
            14'd 2273: out = 12'h4A5;
            14'd 2274: out = 12'h4A5;
            14'd 2275: out = 12'h4A5;
            14'd 2276: out = 12'h4A5;
            14'd 2277: out = 12'h4A5;
            14'd 2278: out = 12'h4A5;
            14'd 2279: out = 12'h4A5;
            14'd 2280: out = 12'h4A6;
            14'd 2281: out = 12'h4A6;
            14'd 2282: out = 12'h4A6;
            14'd 2283: out = 12'h4A6;
            14'd 2284: out = 12'h4A6;
            14'd 2285: out = 12'h4A6;
            14'd 2286: out = 12'h4A6;
            14'd 2287: out = 12'h4A6;
            14'd 2288: out = 12'h4A6;
            14'd 2289: out = 12'h4A6;
            14'd 2290: out = 12'h4A6;
            14'd 2291: out = 12'h4A6;
            14'd 2292: out = 12'h4A7;
            14'd 2293: out = 12'h4A7;
            14'd 2294: out = 12'h4A7;
            14'd 2295: out = 12'h4A7;
            14'd 2296: out = 12'h4A7;
            14'd 2297: out = 12'h4A7;
            14'd 2298: out = 12'h4A7;
            14'd 2299: out = 12'h4A7;
            14'd 2300: out = 12'h4A7;
            14'd 2301: out = 12'h4A7;
            14'd 2302: out = 12'h4A7;
            14'd 2303: out = 12'h4A7;
            14'd 2304: out = 12'h4A8;
            14'd 2305: out = 12'h4A8;
            14'd 2306: out = 12'h4A8;
            14'd 2307: out = 12'h4A8;
            14'd 2308: out = 12'h4A8;
            14'd 2309: out = 12'h4A8;
            14'd 2310: out = 12'h4A8;
            14'd 2311: out = 12'h4A8;
            14'd 2312: out = 12'h4A8;
            14'd 2313: out = 12'h4A8;
            14'd 2314: out = 12'h4A8;
            14'd 2315: out = 12'h4A8;
            14'd 2316: out = 12'h4A9;
            14'd 2317: out = 12'h4A9;
            14'd 2318: out = 12'h4A9;
            14'd 2319: out = 12'h4A9;
            14'd 2320: out = 12'h4A9;
            14'd 2321: out = 12'h4A9;
            14'd 2322: out = 12'h4A9;
            14'd 2323: out = 12'h4A9;
            14'd 2324: out = 12'h4A9;
            14'd 2325: out = 12'h4A9;
            14'd 2326: out = 12'h4A9;
            14'd 2327: out = 12'h4AA;
            14'd 2328: out = 12'h4AA;
            14'd 2329: out = 12'h4AA;
            14'd 2330: out = 12'h4AA;
            14'd 2331: out = 12'h4AA;
            14'd 2332: out = 12'h4AA;
            14'd 2333: out = 12'h4AA;
            14'd 2334: out = 12'h4AA;
            14'd 2335: out = 12'h4AA;
            14'd 2336: out = 12'h4AA;
            14'd 2337: out = 12'h4AA;
            14'd 2338: out = 12'h4AA;
            14'd 2339: out = 12'h4AB;
            14'd 2340: out = 12'h4AB;
            14'd 2341: out = 12'h4AB;
            14'd 2342: out = 12'h4AB;
            14'd 2343: out = 12'h4AB;
            14'd 2344: out = 12'h4AB;
            14'd 2345: out = 12'h4AB;
            14'd 2346: out = 12'h4AB;
            14'd 2347: out = 12'h4AB;
            14'd 2348: out = 12'h4AB;
            14'd 2349: out = 12'h4AB;
            14'd 2350: out = 12'h4AB;
            14'd 2351: out = 12'h4AC;
            14'd 2352: out = 12'h4AC;
            14'd 2353: out = 12'h4AC;
            14'd 2354: out = 12'h4AC;
            14'd 2355: out = 12'h4AC;
            14'd 2356: out = 12'h4AC;
            14'd 2357: out = 12'h4AC;
            14'd 2358: out = 12'h4AC;
            14'd 2359: out = 12'h4AC;
            14'd 2360: out = 12'h4AC;
            14'd 2361: out = 12'h4AC;
            14'd 2362: out = 12'h4AC;
            14'd 2363: out = 12'h4AD;
            14'd 2364: out = 12'h4AD;
            14'd 2365: out = 12'h4AD;
            14'd 2366: out = 12'h4AD;
            14'd 2367: out = 12'h4AD;
            14'd 2368: out = 12'h4AD;
            14'd 2369: out = 12'h4AD;
            14'd 2370: out = 12'h4AD;
            14'd 2371: out = 12'h4AD;
            14'd 2372: out = 12'h4AD;
            14'd 2373: out = 12'h4AD;
            14'd 2374: out = 12'h4AE;
            14'd 2375: out = 12'h4AE;
            14'd 2376: out = 12'h4AE;
            14'd 2377: out = 12'h4AE;
            14'd 2378: out = 12'h4AE;
            14'd 2379: out = 12'h4AE;
            14'd 2380: out = 12'h4AE;
            14'd 2381: out = 12'h4AE;
            14'd 2382: out = 12'h4AE;
            14'd 2383: out = 12'h4AE;
            14'd 2384: out = 12'h4AE;
            14'd 2385: out = 12'h4AE;
            14'd 2386: out = 12'h4AF;
            14'd 2387: out = 12'h4AF;
            14'd 2388: out = 12'h4AF;
            14'd 2389: out = 12'h4AF;
            14'd 2390: out = 12'h4AF;
            14'd 2391: out = 12'h4AF;
            14'd 2392: out = 12'h4AF;
            14'd 2393: out = 12'h4AF;
            14'd 2394: out = 12'h4AF;
            14'd 2395: out = 12'h4AF;
            14'd 2396: out = 12'h4AF;
            14'd 2397: out = 12'h4AF;
            14'd 2398: out = 12'h4B0;
            14'd 2399: out = 12'h4B0;
            14'd 2400: out = 12'h4B0;
            14'd 2401: out = 12'h4B0;
            14'd 2402: out = 12'h4B0;
            14'd 2403: out = 12'h4B0;
            14'd 2404: out = 12'h4B0;
            14'd 2405: out = 12'h4B0;
            14'd 2406: out = 12'h4B0;
            14'd 2407: out = 12'h4B0;
            14'd 2408: out = 12'h4B0;
            14'd 2409: out = 12'h4B1;
            14'd 2410: out = 12'h4B1;
            14'd 2411: out = 12'h4B1;
            14'd 2412: out = 12'h4B1;
            14'd 2413: out = 12'h4B1;
            14'd 2414: out = 12'h4B1;
            14'd 2415: out = 12'h4B1;
            14'd 2416: out = 12'h4B1;
            14'd 2417: out = 12'h4B1;
            14'd 2418: out = 12'h4B1;
            14'd 2419: out = 12'h4B1;
            14'd 2420: out = 12'h4B1;
            14'd 2421: out = 12'h4B2;
            14'd 2422: out = 12'h4B2;
            14'd 2423: out = 12'h4B2;
            14'd 2424: out = 12'h4B2;
            14'd 2425: out = 12'h4B2;
            14'd 2426: out = 12'h4B2;
            14'd 2427: out = 12'h4B2;
            14'd 2428: out = 12'h4B2;
            14'd 2429: out = 12'h4B2;
            14'd 2430: out = 12'h4B2;
            14'd 2431: out = 12'h4B2;
            14'd 2432: out = 12'h4B2;
            14'd 2433: out = 12'h4B3;
            14'd 2434: out = 12'h4B3;
            14'd 2435: out = 12'h4B3;
            14'd 2436: out = 12'h4B3;
            14'd 2437: out = 12'h4B3;
            14'd 2438: out = 12'h4B3;
            14'd 2439: out = 12'h4B3;
            14'd 2440: out = 12'h4B3;
            14'd 2441: out = 12'h4B3;
            14'd 2442: out = 12'h4B3;
            14'd 2443: out = 12'h4B3;
            14'd 2444: out = 12'h4B4;
            14'd 2445: out = 12'h4B4;
            14'd 2446: out = 12'h4B4;
            14'd 2447: out = 12'h4B4;
            14'd 2448: out = 12'h4B4;
            14'd 2449: out = 12'h4B4;
            14'd 2450: out = 12'h4B4;
            14'd 2451: out = 12'h4B4;
            14'd 2452: out = 12'h4B4;
            14'd 2453: out = 12'h4B4;
            14'd 2454: out = 12'h4B4;
            14'd 2455: out = 12'h4B4;
            14'd 2456: out = 12'h4B5;
            14'd 2457: out = 12'h4B5;
            14'd 2458: out = 12'h4B5;
            14'd 2459: out = 12'h4B5;
            14'd 2460: out = 12'h4B5;
            14'd 2461: out = 12'h4B5;
            14'd 2462: out = 12'h4B5;
            14'd 2463: out = 12'h4B5;
            14'd 2464: out = 12'h4B5;
            14'd 2465: out = 12'h4B5;
            14'd 2466: out = 12'h4B5;
            14'd 2467: out = 12'h4B6;
            14'd 2468: out = 12'h4B6;
            14'd 2469: out = 12'h4B6;
            14'd 2470: out = 12'h4B6;
            14'd 2471: out = 12'h4B6;
            14'd 2472: out = 12'h4B6;
            14'd 2473: out = 12'h4B6;
            14'd 2474: out = 12'h4B6;
            14'd 2475: out = 12'h4B6;
            14'd 2476: out = 12'h4B6;
            14'd 2477: out = 12'h4B6;
            14'd 2478: out = 12'h4B6;
            14'd 2479: out = 12'h4B7;
            14'd 2480: out = 12'h4B7;
            14'd 2481: out = 12'h4B7;
            14'd 2482: out = 12'h4B7;
            14'd 2483: out = 12'h4B7;
            14'd 2484: out = 12'h4B7;
            14'd 2485: out = 12'h4B7;
            14'd 2486: out = 12'h4B7;
            14'd 2487: out = 12'h4B7;
            14'd 2488: out = 12'h4B7;
            14'd 2489: out = 12'h4B7;
            14'd 2490: out = 12'h4B8;
            14'd 2491: out = 12'h4B8;
            14'd 2492: out = 12'h4B8;
            14'd 2493: out = 12'h4B8;
            14'd 2494: out = 12'h4B8;
            14'd 2495: out = 12'h4B8;
            14'd 2496: out = 12'h4B8;
            14'd 2497: out = 12'h4B8;
            14'd 2498: out = 12'h4B8;
            14'd 2499: out = 12'h4B8;
            14'd 2500: out = 12'h4B8;
            14'd 2501: out = 12'h4B8;
            14'd 2502: out = 12'h4B9;
            14'd 2503: out = 12'h4B9;
            14'd 2504: out = 12'h4B9;
            14'd 2505: out = 12'h4B9;
            14'd 2506: out = 12'h4B9;
            14'd 2507: out = 12'h4B9;
            14'd 2508: out = 12'h4B9;
            14'd 2509: out = 12'h4B9;
            14'd 2510: out = 12'h4B9;
            14'd 2511: out = 12'h4B9;
            14'd 2512: out = 12'h4B9;
            14'd 2513: out = 12'h4BA;
            14'd 2514: out = 12'h4BA;
            14'd 2515: out = 12'h4BA;
            14'd 2516: out = 12'h4BA;
            14'd 2517: out = 12'h4BA;
            14'd 2518: out = 12'h4BA;
            14'd 2519: out = 12'h4BA;
            14'd 2520: out = 12'h4BA;
            14'd 2521: out = 12'h4BA;
            14'd 2522: out = 12'h4BA;
            14'd 2523: out = 12'h4BA;
            14'd 2524: out = 12'h4BA;
            14'd 2525: out = 12'h4BB;
            14'd 2526: out = 12'h4BB;
            14'd 2527: out = 12'h4BB;
            14'd 2528: out = 12'h4BB;
            14'd 2529: out = 12'h4BB;
            14'd 2530: out = 12'h4BB;
            14'd 2531: out = 12'h4BB;
            14'd 2532: out = 12'h4BB;
            14'd 2533: out = 12'h4BB;
            14'd 2534: out = 12'h4BB;
            14'd 2535: out = 12'h4BB;
            14'd 2536: out = 12'h4BC;
            14'd 2537: out = 12'h4BC;
            14'd 2538: out = 12'h4BC;
            14'd 2539: out = 12'h4BC;
            14'd 2540: out = 12'h4BC;
            14'd 2541: out = 12'h4BC;
            14'd 2542: out = 12'h4BC;
            14'd 2543: out = 12'h4BC;
            14'd 2544: out = 12'h4BC;
            14'd 2545: out = 12'h4BC;
            14'd 2546: out = 12'h4BC;
            14'd 2547: out = 12'h4BC;
            14'd 2548: out = 12'h4BD;
            14'd 2549: out = 12'h4BD;
            14'd 2550: out = 12'h4BD;
            14'd 2551: out = 12'h4BD;
            14'd 2552: out = 12'h4BD;
            14'd 2553: out = 12'h4BD;
            14'd 2554: out = 12'h4BD;
            14'd 2555: out = 12'h4BD;
            14'd 2556: out = 12'h4BD;
            14'd 2557: out = 12'h4BD;
            14'd 2558: out = 12'h4BD;
            14'd 2559: out = 12'h4BE;
            14'd 2560: out = 12'h4BE;
            14'd 2561: out = 12'h4BE;
            14'd 2562: out = 12'h4BE;
            14'd 2563: out = 12'h4BE;
            14'd 2564: out = 12'h4BE;
            14'd 2565: out = 12'h4BE;
            14'd 2566: out = 12'h4BE;
            14'd 2567: out = 12'h4BE;
            14'd 2568: out = 12'h4BE;
            14'd 2569: out = 12'h4BE;
            14'd 2570: out = 12'h4BF;
            14'd 2571: out = 12'h4BF;
            14'd 2572: out = 12'h4BF;
            14'd 2573: out = 12'h4BF;
            14'd 2574: out = 12'h4BF;
            14'd 2575: out = 12'h4BF;
            14'd 2576: out = 12'h4BF;
            14'd 2577: out = 12'h4BF;
            14'd 2578: out = 12'h4BF;
            14'd 2579: out = 12'h4BF;
            14'd 2580: out = 12'h4BF;
            14'd 2581: out = 12'h4BF;
            14'd 2582: out = 12'h4C0;
            14'd 2583: out = 12'h4C0;
            14'd 2584: out = 12'h4C0;
            14'd 2585: out = 12'h4C0;
            14'd 2586: out = 12'h4C0;
            14'd 2587: out = 12'h4C0;
            14'd 2588: out = 12'h4C0;
            14'd 2589: out = 12'h4C0;
            14'd 2590: out = 12'h4C0;
            14'd 2591: out = 12'h4C0;
            14'd 2592: out = 12'h4C0;
            14'd 2593: out = 12'h4C1;
            14'd 2594: out = 12'h4C1;
            14'd 2595: out = 12'h4C1;
            14'd 2596: out = 12'h4C1;
            14'd 2597: out = 12'h4C1;
            14'd 2598: out = 12'h4C1;
            14'd 2599: out = 12'h4C1;
            14'd 2600: out = 12'h4C1;
            14'd 2601: out = 12'h4C1;
            14'd 2602: out = 12'h4C1;
            14'd 2603: out = 12'h4C1;
            14'd 2604: out = 12'h4C2;
            14'd 2605: out = 12'h4C2;
            14'd 2606: out = 12'h4C2;
            14'd 2607: out = 12'h4C2;
            14'd 2608: out = 12'h4C2;
            14'd 2609: out = 12'h4C2;
            14'd 2610: out = 12'h4C2;
            14'd 2611: out = 12'h4C2;
            14'd 2612: out = 12'h4C2;
            14'd 2613: out = 12'h4C2;
            14'd 2614: out = 12'h4C2;
            14'd 2615: out = 12'h4C2;
            14'd 2616: out = 12'h4C3;
            14'd 2617: out = 12'h4C3;
            14'd 2618: out = 12'h4C3;
            14'd 2619: out = 12'h4C3;
            14'd 2620: out = 12'h4C3;
            14'd 2621: out = 12'h4C3;
            14'd 2622: out = 12'h4C3;
            14'd 2623: out = 12'h4C3;
            14'd 2624: out = 12'h4C3;
            14'd 2625: out = 12'h4C3;
            14'd 2626: out = 12'h4C3;
            14'd 2627: out = 12'h4C4;
            14'd 2628: out = 12'h4C4;
            14'd 2629: out = 12'h4C4;
            14'd 2630: out = 12'h4C4;
            14'd 2631: out = 12'h4C4;
            14'd 2632: out = 12'h4C4;
            14'd 2633: out = 12'h4C4;
            14'd 2634: out = 12'h4C4;
            14'd 2635: out = 12'h4C4;
            14'd 2636: out = 12'h4C4;
            14'd 2637: out = 12'h4C4;
            14'd 2638: out = 12'h4C5;
            14'd 2639: out = 12'h4C5;
            14'd 2640: out = 12'h4C5;
            14'd 2641: out = 12'h4C5;
            14'd 2642: out = 12'h4C5;
            14'd 2643: out = 12'h4C5;
            14'd 2644: out = 12'h4C5;
            14'd 2645: out = 12'h4C5;
            14'd 2646: out = 12'h4C5;
            14'd 2647: out = 12'h4C5;
            14'd 2648: out = 12'h4C5;
            14'd 2649: out = 12'h4C5;
            14'd 2650: out = 12'h4C6;
            14'd 2651: out = 12'h4C6;
            14'd 2652: out = 12'h4C6;
            14'd 2653: out = 12'h4C6;
            14'd 2654: out = 12'h4C6;
            14'd 2655: out = 12'h4C6;
            14'd 2656: out = 12'h4C6;
            14'd 2657: out = 12'h4C6;
            14'd 2658: out = 12'h4C6;
            14'd 2659: out = 12'h4C6;
            14'd 2660: out = 12'h4C6;
            14'd 2661: out = 12'h4C7;
            14'd 2662: out = 12'h4C7;
            14'd 2663: out = 12'h4C7;
            14'd 2664: out = 12'h4C7;
            14'd 2665: out = 12'h4C7;
            14'd 2666: out = 12'h4C7;
            14'd 2667: out = 12'h4C7;
            14'd 2668: out = 12'h4C7;
            14'd 2669: out = 12'h4C7;
            14'd 2670: out = 12'h4C7;
            14'd 2671: out = 12'h4C7;
            14'd 2672: out = 12'h4C8;
            14'd 2673: out = 12'h4C8;
            14'd 2674: out = 12'h4C8;
            14'd 2675: out = 12'h4C8;
            14'd 2676: out = 12'h4C8;
            14'd 2677: out = 12'h4C8;
            14'd 2678: out = 12'h4C8;
            14'd 2679: out = 12'h4C8;
            14'd 2680: out = 12'h4C8;
            14'd 2681: out = 12'h4C8;
            14'd 2682: out = 12'h4C8;
            14'd 2683: out = 12'h4C9;
            14'd 2684: out = 12'h4C9;
            14'd 2685: out = 12'h4C9;
            14'd 2686: out = 12'h4C9;
            14'd 2687: out = 12'h4C9;
            14'd 2688: out = 12'h4C9;
            14'd 2689: out = 12'h4C9;
            14'd 2690: out = 12'h4C9;
            14'd 2691: out = 12'h4C9;
            14'd 2692: out = 12'h4C9;
            14'd 2693: out = 12'h4C9;
            14'd 2694: out = 12'h4CA;
            14'd 2695: out = 12'h4CA;
            14'd 2696: out = 12'h4CA;
            14'd 2697: out = 12'h4CA;
            14'd 2698: out = 12'h4CA;
            14'd 2699: out = 12'h4CA;
            14'd 2700: out = 12'h4CA;
            14'd 2701: out = 12'h4CA;
            14'd 2702: out = 12'h4CA;
            14'd 2703: out = 12'h4CA;
            14'd 2704: out = 12'h4CA;
            14'd 2705: out = 12'h4CA;
            14'd 2706: out = 12'h4CB;
            14'd 2707: out = 12'h4CB;
            14'd 2708: out = 12'h4CB;
            14'd 2709: out = 12'h4CB;
            14'd 2710: out = 12'h4CB;
            14'd 2711: out = 12'h4CB;
            14'd 2712: out = 12'h4CB;
            14'd 2713: out = 12'h4CB;
            14'd 2714: out = 12'h4CB;
            14'd 2715: out = 12'h4CB;
            14'd 2716: out = 12'h4CB;
            14'd 2717: out = 12'h4CC;
            14'd 2718: out = 12'h4CC;
            14'd 2719: out = 12'h4CC;
            14'd 2720: out = 12'h4CC;
            14'd 2721: out = 12'h4CC;
            14'd 2722: out = 12'h4CC;
            14'd 2723: out = 12'h4CC;
            14'd 2724: out = 12'h4CC;
            14'd 2725: out = 12'h4CC;
            14'd 2726: out = 12'h4CC;
            14'd 2727: out = 12'h4CC;
            14'd 2728: out = 12'h4CD;
            14'd 2729: out = 12'h4CD;
            14'd 2730: out = 12'h4CD;
            14'd 2731: out = 12'h4CD;
            14'd 2732: out = 12'h4CD;
            14'd 2733: out = 12'h4CD;
            14'd 2734: out = 12'h4CD;
            14'd 2735: out = 12'h4CD;
            14'd 2736: out = 12'h4CD;
            14'd 2737: out = 12'h4CD;
            14'd 2738: out = 12'h4CD;
            14'd 2739: out = 12'h4CE;
            14'd 2740: out = 12'h4CE;
            14'd 2741: out = 12'h4CE;
            14'd 2742: out = 12'h4CE;
            14'd 2743: out = 12'h4CE;
            14'd 2744: out = 12'h4CE;
            14'd 2745: out = 12'h4CE;
            14'd 2746: out = 12'h4CE;
            14'd 2747: out = 12'h4CE;
            14'd 2748: out = 12'h4CE;
            14'd 2749: out = 12'h4CE;
            14'd 2750: out = 12'h4CF;
            14'd 2751: out = 12'h4CF;
            14'd 2752: out = 12'h4CF;
            14'd 2753: out = 12'h4CF;
            14'd 2754: out = 12'h4CF;
            14'd 2755: out = 12'h4CF;
            14'd 2756: out = 12'h4CF;
            14'd 2757: out = 12'h4CF;
            14'd 2758: out = 12'h4CF;
            14'd 2759: out = 12'h4CF;
            14'd 2760: out = 12'h4CF;
            14'd 2761: out = 12'h4D0;
            14'd 2762: out = 12'h4D0;
            14'd 2763: out = 12'h4D0;
            14'd 2764: out = 12'h4D0;
            14'd 2765: out = 12'h4D0;
            14'd 2766: out = 12'h4D0;
            14'd 2767: out = 12'h4D0;
            14'd 2768: out = 12'h4D0;
            14'd 2769: out = 12'h4D0;
            14'd 2770: out = 12'h4D0;
            14'd 2771: out = 12'h4D0;
            14'd 2772: out = 12'h4D1;
            14'd 2773: out = 12'h4D1;
            14'd 2774: out = 12'h4D1;
            14'd 2775: out = 12'h4D1;
            14'd 2776: out = 12'h4D1;
            14'd 2777: out = 12'h4D1;
            14'd 2778: out = 12'h4D1;
            14'd 2779: out = 12'h4D1;
            14'd 2780: out = 12'h4D1;
            14'd 2781: out = 12'h4D1;
            14'd 2782: out = 12'h4D1;
            14'd 2783: out = 12'h4D2;
            14'd 2784: out = 12'h4D2;
            14'd 2785: out = 12'h4D2;
            14'd 2786: out = 12'h4D2;
            14'd 2787: out = 12'h4D2;
            14'd 2788: out = 12'h4D2;
            14'd 2789: out = 12'h4D2;
            14'd 2790: out = 12'h4D2;
            14'd 2791: out = 12'h4D2;
            14'd 2792: out = 12'h4D2;
            14'd 2793: out = 12'h4D2;
            14'd 2794: out = 12'h4D3;
            14'd 2795: out = 12'h4D3;
            14'd 2796: out = 12'h4D3;
            14'd 2797: out = 12'h4D3;
            14'd 2798: out = 12'h4D3;
            14'd 2799: out = 12'h4D3;
            14'd 2800: out = 12'h4D3;
            14'd 2801: out = 12'h4D3;
            14'd 2802: out = 12'h4D3;
            14'd 2803: out = 12'h4D3;
            14'd 2804: out = 12'h4D3;
            14'd 2805: out = 12'h4D4;
            14'd 2806: out = 12'h4D4;
            14'd 2807: out = 12'h4D4;
            14'd 2808: out = 12'h4D4;
            14'd 2809: out = 12'h4D4;
            14'd 2810: out = 12'h4D4;
            14'd 2811: out = 12'h4D4;
            14'd 2812: out = 12'h4D4;
            14'd 2813: out = 12'h4D4;
            14'd 2814: out = 12'h4D4;
            14'd 2815: out = 12'h4D4;
            14'd 2816: out = 12'h4D5;
            14'd 2817: out = 12'h4D5;
            14'd 2818: out = 12'h4D5;
            14'd 2819: out = 12'h4D5;
            14'd 2820: out = 12'h4D5;
            14'd 2821: out = 12'h4D5;
            14'd 2822: out = 12'h4D5;
            14'd 2823: out = 12'h4D5;
            14'd 2824: out = 12'h4D5;
            14'd 2825: out = 12'h4D5;
            14'd 2826: out = 12'h4D5;
            14'd 2827: out = 12'h4D6;
            14'd 2828: out = 12'h4D6;
            14'd 2829: out = 12'h4D6;
            14'd 2830: out = 12'h4D6;
            14'd 2831: out = 12'h4D6;
            14'd 2832: out = 12'h4D6;
            14'd 2833: out = 12'h4D6;
            14'd 2834: out = 12'h4D6;
            14'd 2835: out = 12'h4D6;
            14'd 2836: out = 12'h4D6;
            14'd 2837: out = 12'h4D6;
            14'd 2838: out = 12'h4D7;
            14'd 2839: out = 12'h4D7;
            14'd 2840: out = 12'h4D7;
            14'd 2841: out = 12'h4D7;
            14'd 2842: out = 12'h4D7;
            14'd 2843: out = 12'h4D7;
            14'd 2844: out = 12'h4D7;
            14'd 2845: out = 12'h4D7;
            14'd 2846: out = 12'h4D7;
            14'd 2847: out = 12'h4D7;
            14'd 2848: out = 12'h4D7;
            14'd 2849: out = 12'h4D8;
            14'd 2850: out = 12'h4D8;
            14'd 2851: out = 12'h4D8;
            14'd 2852: out = 12'h4D8;
            14'd 2853: out = 12'h4D8;
            14'd 2854: out = 12'h4D8;
            14'd 2855: out = 12'h4D8;
            14'd 2856: out = 12'h4D8;
            14'd 2857: out = 12'h4D8;
            14'd 2858: out = 12'h4D8;
            14'd 2859: out = 12'h4D8;
            14'd 2860: out = 12'h4D9;
            14'd 2861: out = 12'h4D9;
            14'd 2862: out = 12'h4D9;
            14'd 2863: out = 12'h4D9;
            14'd 2864: out = 12'h4D9;
            14'd 2865: out = 12'h4D9;
            14'd 2866: out = 12'h4D9;
            14'd 2867: out = 12'h4D9;
            14'd 2868: out = 12'h4D9;
            14'd 2869: out = 12'h4D9;
            14'd 2870: out = 12'h4D9;
            14'd 2871: out = 12'h4DA;
            14'd 2872: out = 12'h4DA;
            14'd 2873: out = 12'h4DA;
            14'd 2874: out = 12'h4DA;
            14'd 2875: out = 12'h4DA;
            14'd 2876: out = 12'h4DA;
            14'd 2877: out = 12'h4DA;
            14'd 2878: out = 12'h4DA;
            14'd 2879: out = 12'h4DA;
            14'd 2880: out = 12'h4DA;
            14'd 2881: out = 12'h4DA;
            14'd 2882: out = 12'h4DB;
            14'd 2883: out = 12'h4DB;
            14'd 2884: out = 12'h4DB;
            14'd 2885: out = 12'h4DB;
            14'd 2886: out = 12'h4DB;
            14'd 2887: out = 12'h4DB;
            14'd 2888: out = 12'h4DB;
            14'd 2889: out = 12'h4DB;
            14'd 2890: out = 12'h4DB;
            14'd 2891: out = 12'h4DB;
            14'd 2892: out = 12'h4DB;
            14'd 2893: out = 12'h4DC;
            14'd 2894: out = 12'h4DC;
            14'd 2895: out = 12'h4DC;
            14'd 2896: out = 12'h4DC;
            14'd 2897: out = 12'h4DC;
            14'd 2898: out = 12'h4DC;
            14'd 2899: out = 12'h4DC;
            14'd 2900: out = 12'h4DC;
            14'd 2901: out = 12'h4DC;
            14'd 2902: out = 12'h4DC;
            14'd 2903: out = 12'h4DD;
            14'd 2904: out = 12'h4DD;
            14'd 2905: out = 12'h4DD;
            14'd 2906: out = 12'h4DD;
            14'd 2907: out = 12'h4DD;
            14'd 2908: out = 12'h4DD;
            14'd 2909: out = 12'h4DD;
            14'd 2910: out = 12'h4DD;
            14'd 2911: out = 12'h4DD;
            14'd 2912: out = 12'h4DD;
            14'd 2913: out = 12'h4DD;
            14'd 2914: out = 12'h4DE;
            14'd 2915: out = 12'h4DE;
            14'd 2916: out = 12'h4DE;
            14'd 2917: out = 12'h4DE;
            14'd 2918: out = 12'h4DE;
            14'd 2919: out = 12'h4DE;
            14'd 2920: out = 12'h4DE;
            14'd 2921: out = 12'h4DE;
            14'd 2922: out = 12'h4DE;
            14'd 2923: out = 12'h4DE;
            14'd 2924: out = 12'h4DE;
            14'd 2925: out = 12'h4DF;
            14'd 2926: out = 12'h4DF;
            14'd 2927: out = 12'h4DF;
            14'd 2928: out = 12'h4DF;
            14'd 2929: out = 12'h4DF;
            14'd 2930: out = 12'h4DF;
            14'd 2931: out = 12'h4DF;
            14'd 2932: out = 12'h4DF;
            14'd 2933: out = 12'h4DF;
            14'd 2934: out = 12'h4DF;
            14'd 2935: out = 12'h4DF;
            14'd 2936: out = 12'h4E0;
            14'd 2937: out = 12'h4E0;
            14'd 2938: out = 12'h4E0;
            14'd 2939: out = 12'h4E0;
            14'd 2940: out = 12'h4E0;
            14'd 2941: out = 12'h4E0;
            14'd 2942: out = 12'h4E0;
            14'd 2943: out = 12'h4E0;
            14'd 2944: out = 12'h4E0;
            14'd 2945: out = 12'h4E0;
            14'd 2946: out = 12'h4E0;
            14'd 2947: out = 12'h4E1;
            14'd 2948: out = 12'h4E1;
            14'd 2949: out = 12'h4E1;
            14'd 2950: out = 12'h4E1;
            14'd 2951: out = 12'h4E1;
            14'd 2952: out = 12'h4E1;
            14'd 2953: out = 12'h4E1;
            14'd 2954: out = 12'h4E1;
            14'd 2955: out = 12'h4E1;
            14'd 2956: out = 12'h4E1;
            14'd 2957: out = 12'h4E2;
            14'd 2958: out = 12'h4E2;
            14'd 2959: out = 12'h4E2;
            14'd 2960: out = 12'h4E2;
            14'd 2961: out = 12'h4E2;
            14'd 2962: out = 12'h4E2;
            14'd 2963: out = 12'h4E2;
            14'd 2964: out = 12'h4E2;
            14'd 2965: out = 12'h4E2;
            14'd 2966: out = 12'h4E2;
            14'd 2967: out = 12'h4E2;
            14'd 2968: out = 12'h4E3;
            14'd 2969: out = 12'h4E3;
            14'd 2970: out = 12'h4E3;
            14'd 2971: out = 12'h4E3;
            14'd 2972: out = 12'h4E3;
            14'd 2973: out = 12'h4E3;
            14'd 2974: out = 12'h4E3;
            14'd 2975: out = 12'h4E3;
            14'd 2976: out = 12'h4E3;
            14'd 2977: out = 12'h4E3;
            14'd 2978: out = 12'h4E3;
            14'd 2979: out = 12'h4E4;
            14'd 2980: out = 12'h4E4;
            14'd 2981: out = 12'h4E4;
            14'd 2982: out = 12'h4E4;
            14'd 2983: out = 12'h4E4;
            14'd 2984: out = 12'h4E4;
            14'd 2985: out = 12'h4E4;
            14'd 2986: out = 12'h4E4;
            14'd 2987: out = 12'h4E4;
            14'd 2988: out = 12'h4E4;
            14'd 2989: out = 12'h4E4;
            14'd 2990: out = 12'h4E5;
            14'd 2991: out = 12'h4E5;
            14'd 2992: out = 12'h4E5;
            14'd 2993: out = 12'h4E5;
            14'd 2994: out = 12'h4E5;
            14'd 2995: out = 12'h4E5;
            14'd 2996: out = 12'h4E5;
            14'd 2997: out = 12'h4E5;
            14'd 2998: out = 12'h4E5;
            14'd 2999: out = 12'h4E5;
            14'd 3000: out = 12'h4E6;
            14'd 3001: out = 12'h4E6;
            14'd 3002: out = 12'h4E6;
            14'd 3003: out = 12'h4E6;
            14'd 3004: out = 12'h4E6;
            14'd 3005: out = 12'h4E6;
            14'd 3006: out = 12'h4E6;
            14'd 3007: out = 12'h4E6;
            14'd 3008: out = 12'h4E6;
            14'd 3009: out = 12'h4E6;
            14'd 3010: out = 12'h4E6;
            14'd 3011: out = 12'h4E7;
            14'd 3012: out = 12'h4E7;
            14'd 3013: out = 12'h4E7;
            14'd 3014: out = 12'h4E7;
            14'd 3015: out = 12'h4E7;
            14'd 3016: out = 12'h4E7;
            14'd 3017: out = 12'h4E7;
            14'd 3018: out = 12'h4E7;
            14'd 3019: out = 12'h4E7;
            14'd 3020: out = 12'h4E7;
            14'd 3021: out = 12'h4E7;
            14'd 3022: out = 12'h4E8;
            14'd 3023: out = 12'h4E8;
            14'd 3024: out = 12'h4E8;
            14'd 3025: out = 12'h4E8;
            14'd 3026: out = 12'h4E8;
            14'd 3027: out = 12'h4E8;
            14'd 3028: out = 12'h4E8;
            14'd 3029: out = 12'h4E8;
            14'd 3030: out = 12'h4E8;
            14'd 3031: out = 12'h4E8;
            14'd 3032: out = 12'h4E9;
            14'd 3033: out = 12'h4E9;
            14'd 3034: out = 12'h4E9;
            14'd 3035: out = 12'h4E9;
            14'd 3036: out = 12'h4E9;
            14'd 3037: out = 12'h4E9;
            14'd 3038: out = 12'h4E9;
            14'd 3039: out = 12'h4E9;
            14'd 3040: out = 12'h4E9;
            14'd 3041: out = 12'h4E9;
            14'd 3042: out = 12'h4E9;
            14'd 3043: out = 12'h4EA;
            14'd 3044: out = 12'h4EA;
            14'd 3045: out = 12'h4EA;
            14'd 3046: out = 12'h4EA;
            14'd 3047: out = 12'h4EA;
            14'd 3048: out = 12'h4EA;
            14'd 3049: out = 12'h4EA;
            14'd 3050: out = 12'h4EA;
            14'd 3051: out = 12'h4EA;
            14'd 3052: out = 12'h4EA;
            14'd 3053: out = 12'h4EB;
            14'd 3054: out = 12'h4EB;
            14'd 3055: out = 12'h4EB;
            14'd 3056: out = 12'h4EB;
            14'd 3057: out = 12'h4EB;
            14'd 3058: out = 12'h4EB;
            14'd 3059: out = 12'h4EB;
            14'd 3060: out = 12'h4EB;
            14'd 3061: out = 12'h4EB;
            14'd 3062: out = 12'h4EB;
            14'd 3063: out = 12'h4EB;
            14'd 3064: out = 12'h4EC;
            14'd 3065: out = 12'h4EC;
            14'd 3066: out = 12'h4EC;
            14'd 3067: out = 12'h4EC;
            14'd 3068: out = 12'h4EC;
            14'd 3069: out = 12'h4EC;
            14'd 3070: out = 12'h4EC;
            14'd 3071: out = 12'h4EC;
            14'd 3072: out = 12'h4EC;
            14'd 3073: out = 12'h4EC;
            14'd 3074: out = 12'h4EC;
            14'd 3075: out = 12'h4ED;
            14'd 3076: out = 12'h4ED;
            14'd 3077: out = 12'h4ED;
            14'd 3078: out = 12'h4ED;
            14'd 3079: out = 12'h4ED;
            14'd 3080: out = 12'h4ED;
            14'd 3081: out = 12'h4ED;
            14'd 3082: out = 12'h4ED;
            14'd 3083: out = 12'h4ED;
            14'd 3084: out = 12'h4ED;
            14'd 3085: out = 12'h4EE;
            14'd 3086: out = 12'h4EE;
            14'd 3087: out = 12'h4EE;
            14'd 3088: out = 12'h4EE;
            14'd 3089: out = 12'h4EE;
            14'd 3090: out = 12'h4EE;
            14'd 3091: out = 12'h4EE;
            14'd 3092: out = 12'h4EE;
            14'd 3093: out = 12'h4EE;
            14'd 3094: out = 12'h4EE;
            14'd 3095: out = 12'h4EE;
            14'd 3096: out = 12'h4EF;
            14'd 3097: out = 12'h4EF;
            14'd 3098: out = 12'h4EF;
            14'd 3099: out = 12'h4EF;
            14'd 3100: out = 12'h4EF;
            14'd 3101: out = 12'h4EF;
            14'd 3102: out = 12'h4EF;
            14'd 3103: out = 12'h4EF;
            14'd 3104: out = 12'h4EF;
            14'd 3105: out = 12'h4EF;
            14'd 3106: out = 12'h4F0;
            14'd 3107: out = 12'h4F0;
            14'd 3108: out = 12'h4F0;
            14'd 3109: out = 12'h4F0;
            14'd 3110: out = 12'h4F0;
            14'd 3111: out = 12'h4F0;
            14'd 3112: out = 12'h4F0;
            14'd 3113: out = 12'h4F0;
            14'd 3114: out = 12'h4F0;
            14'd 3115: out = 12'h4F0;
            14'd 3116: out = 12'h4F0;
            14'd 3117: out = 12'h4F1;
            14'd 3118: out = 12'h4F1;
            14'd 3119: out = 12'h4F1;
            14'd 3120: out = 12'h4F1;
            14'd 3121: out = 12'h4F1;
            14'd 3122: out = 12'h4F1;
            14'd 3123: out = 12'h4F1;
            14'd 3124: out = 12'h4F1;
            14'd 3125: out = 12'h4F1;
            14'd 3126: out = 12'h4F1;
            14'd 3127: out = 12'h4F2;
            14'd 3128: out = 12'h4F2;
            14'd 3129: out = 12'h4F2;
            14'd 3130: out = 12'h4F2;
            14'd 3131: out = 12'h4F2;
            14'd 3132: out = 12'h4F2;
            14'd 3133: out = 12'h4F2;
            14'd 3134: out = 12'h4F2;
            14'd 3135: out = 12'h4F2;
            14'd 3136: out = 12'h4F2;
            14'd 3137: out = 12'h4F2;
            14'd 3138: out = 12'h4F3;
            14'd 3139: out = 12'h4F3;
            14'd 3140: out = 12'h4F3;
            14'd 3141: out = 12'h4F3;
            14'd 3142: out = 12'h4F3;
            14'd 3143: out = 12'h4F3;
            14'd 3144: out = 12'h4F3;
            14'd 3145: out = 12'h4F3;
            14'd 3146: out = 12'h4F3;
            14'd 3147: out = 12'h4F3;
            14'd 3148: out = 12'h4F4;
            14'd 3149: out = 12'h4F4;
            14'd 3150: out = 12'h4F4;
            14'd 3151: out = 12'h4F4;
            14'd 3152: out = 12'h4F4;
            14'd 3153: out = 12'h4F4;
            14'd 3154: out = 12'h4F4;
            14'd 3155: out = 12'h4F4;
            14'd 3156: out = 12'h4F4;
            14'd 3157: out = 12'h4F4;
            14'd 3158: out = 12'h4F5;
            14'd 3159: out = 12'h4F5;
            14'd 3160: out = 12'h4F5;
            14'd 3161: out = 12'h4F5;
            14'd 3162: out = 12'h4F5;
            14'd 3163: out = 12'h4F5;
            14'd 3164: out = 12'h4F5;
            14'd 3165: out = 12'h4F5;
            14'd 3166: out = 12'h4F5;
            14'd 3167: out = 12'h4F5;
            14'd 3168: out = 12'h4F5;
            14'd 3169: out = 12'h4F6;
            14'd 3170: out = 12'h4F6;
            14'd 3171: out = 12'h4F6;
            14'd 3172: out = 12'h4F6;
            14'd 3173: out = 12'h4F6;
            14'd 3174: out = 12'h4F6;
            14'd 3175: out = 12'h4F6;
            14'd 3176: out = 12'h4F6;
            14'd 3177: out = 12'h4F6;
            14'd 3178: out = 12'h4F6;
            14'd 3179: out = 12'h4F7;
            14'd 3180: out = 12'h4F7;
            14'd 3181: out = 12'h4F7;
            14'd 3182: out = 12'h4F7;
            14'd 3183: out = 12'h4F7;
            14'd 3184: out = 12'h4F7;
            14'd 3185: out = 12'h4F7;
            14'd 3186: out = 12'h4F7;
            14'd 3187: out = 12'h4F7;
            14'd 3188: out = 12'h4F7;
            14'd 3189: out = 12'h4F7;
            14'd 3190: out = 12'h4F8;
            14'd 3191: out = 12'h4F8;
            14'd 3192: out = 12'h4F8;
            14'd 3193: out = 12'h4F8;
            14'd 3194: out = 12'h4F8;
            14'd 3195: out = 12'h4F8;
            14'd 3196: out = 12'h4F8;
            14'd 3197: out = 12'h4F8;
            14'd 3198: out = 12'h4F8;
            14'd 3199: out = 12'h4F8;
            14'd 3200: out = 12'h4F9;
            14'd 3201: out = 12'h4F9;
            14'd 3202: out = 12'h4F9;
            14'd 3203: out = 12'h4F9;
            14'd 3204: out = 12'h4F9;
            14'd 3205: out = 12'h4F9;
            14'd 3206: out = 12'h4F9;
            14'd 3207: out = 12'h4F9;
            14'd 3208: out = 12'h4F9;
            14'd 3209: out = 12'h4F9;
            14'd 3210: out = 12'h4FA;
            14'd 3211: out = 12'h4FA;
            14'd 3212: out = 12'h4FA;
            14'd 3213: out = 12'h4FA;
            14'd 3214: out = 12'h4FA;
            14'd 3215: out = 12'h4FA;
            14'd 3216: out = 12'h4FA;
            14'd 3217: out = 12'h4FA;
            14'd 3218: out = 12'h4FA;
            14'd 3219: out = 12'h4FA;
            14'd 3220: out = 12'h4FA;
            14'd 3221: out = 12'h4FB;
            14'd 3222: out = 12'h4FB;
            14'd 3223: out = 12'h4FB;
            14'd 3224: out = 12'h4FB;
            14'd 3225: out = 12'h4FB;
            14'd 3226: out = 12'h4FB;
            14'd 3227: out = 12'h4FB;
            14'd 3228: out = 12'h4FB;
            14'd 3229: out = 12'h4FB;
            14'd 3230: out = 12'h4FB;
            14'd 3231: out = 12'h4FC;
            14'd 3232: out = 12'h4FC;
            14'd 3233: out = 12'h4FC;
            14'd 3234: out = 12'h4FC;
            14'd 3235: out = 12'h4FC;
            14'd 3236: out = 12'h4FC;
            14'd 3237: out = 12'h4FC;
            14'd 3238: out = 12'h4FC;
            14'd 3239: out = 12'h4FC;
            14'd 3240: out = 12'h4FC;
            14'd 3241: out = 12'h4FD;
            14'd 3242: out = 12'h4FD;
            14'd 3243: out = 12'h4FD;
            14'd 3244: out = 12'h4FD;
            14'd 3245: out = 12'h4FD;
            14'd 3246: out = 12'h4FD;
            14'd 3247: out = 12'h4FD;
            14'd 3248: out = 12'h4FD;
            14'd 3249: out = 12'h4FD;
            14'd 3250: out = 12'h4FD;
            14'd 3251: out = 12'h4FD;
            14'd 3252: out = 12'h4FE;
            14'd 3253: out = 12'h4FE;
            14'd 3254: out = 12'h4FE;
            14'd 3255: out = 12'h4FE;
            14'd 3256: out = 12'h4FE;
            14'd 3257: out = 12'h4FE;
            14'd 3258: out = 12'h4FE;
            14'd 3259: out = 12'h4FE;
            14'd 3260: out = 12'h4FE;
            14'd 3261: out = 12'h4FE;
            14'd 3262: out = 12'h4FF;
            14'd 3263: out = 12'h4FF;
            14'd 3264: out = 12'h4FF;
            14'd 3265: out = 12'h4FF;
            14'd 3266: out = 12'h4FF;
            14'd 3267: out = 12'h4FF;
            14'd 3268: out = 12'h4FF;
            14'd 3269: out = 12'h4FF;
            14'd 3270: out = 12'h4FF;
            14'd 3271: out = 12'h4FF;
            14'd 3272: out = 12'h500;
            14'd 3273: out = 12'h500;
            14'd 3274: out = 12'h500;
            14'd 3275: out = 12'h500;
            14'd 3276: out = 12'h500;
            14'd 3277: out = 12'h500;
            14'd 3278: out = 12'h500;
            14'd 3279: out = 12'h500;
            14'd 3280: out = 12'h500;
            14'd 3281: out = 12'h500;
            14'd 3282: out = 12'h501;
            14'd 3283: out = 12'h501;
            14'd 3284: out = 12'h501;
            14'd 3285: out = 12'h501;
            14'd 3286: out = 12'h501;
            14'd 3287: out = 12'h501;
            14'd 3288: out = 12'h501;
            14'd 3289: out = 12'h501;
            14'd 3290: out = 12'h501;
            14'd 3291: out = 12'h501;
            14'd 3292: out = 12'h501;
            14'd 3293: out = 12'h502;
            14'd 3294: out = 12'h502;
            14'd 3295: out = 12'h502;
            14'd 3296: out = 12'h502;
            14'd 3297: out = 12'h502;
            14'd 3298: out = 12'h502;
            14'd 3299: out = 12'h502;
            14'd 3300: out = 12'h502;
            14'd 3301: out = 12'h502;
            14'd 3302: out = 12'h502;
            14'd 3303: out = 12'h503;
            14'd 3304: out = 12'h503;
            14'd 3305: out = 12'h503;
            14'd 3306: out = 12'h503;
            14'd 3307: out = 12'h503;
            14'd 3308: out = 12'h503;
            14'd 3309: out = 12'h503;
            14'd 3310: out = 12'h503;
            14'd 3311: out = 12'h503;
            14'd 3312: out = 12'h503;
            14'd 3313: out = 12'h504;
            14'd 3314: out = 12'h504;
            14'd 3315: out = 12'h504;
            14'd 3316: out = 12'h504;
            14'd 3317: out = 12'h504;
            14'd 3318: out = 12'h504;
            14'd 3319: out = 12'h504;
            14'd 3320: out = 12'h504;
            14'd 3321: out = 12'h504;
            14'd 3322: out = 12'h504;
            14'd 3323: out = 12'h505;
            14'd 3324: out = 12'h505;
            14'd 3325: out = 12'h505;
            14'd 3326: out = 12'h505;
            14'd 3327: out = 12'h505;
            14'd 3328: out = 12'h505;
            14'd 3329: out = 12'h505;
            14'd 3330: out = 12'h505;
            14'd 3331: out = 12'h505;
            14'd 3332: out = 12'h505;
            14'd 3333: out = 12'h506;
            14'd 3334: out = 12'h506;
            14'd 3335: out = 12'h506;
            14'd 3336: out = 12'h506;
            14'd 3337: out = 12'h506;
            14'd 3338: out = 12'h506;
            14'd 3339: out = 12'h506;
            14'd 3340: out = 12'h506;
            14'd 3341: out = 12'h506;
            14'd 3342: out = 12'h506;
            14'd 3343: out = 12'h506;
            14'd 3344: out = 12'h507;
            14'd 3345: out = 12'h507;
            14'd 3346: out = 12'h507;
            14'd 3347: out = 12'h507;
            14'd 3348: out = 12'h507;
            14'd 3349: out = 12'h507;
            14'd 3350: out = 12'h507;
            14'd 3351: out = 12'h507;
            14'd 3352: out = 12'h507;
            14'd 3353: out = 12'h507;
            14'd 3354: out = 12'h508;
            14'd 3355: out = 12'h508;
            14'd 3356: out = 12'h508;
            14'd 3357: out = 12'h508;
            14'd 3358: out = 12'h508;
            14'd 3359: out = 12'h508;
            14'd 3360: out = 12'h508;
            14'd 3361: out = 12'h508;
            14'd 3362: out = 12'h508;
            14'd 3363: out = 12'h508;
            14'd 3364: out = 12'h509;
            14'd 3365: out = 12'h509;
            14'd 3366: out = 12'h509;
            14'd 3367: out = 12'h509;
            14'd 3368: out = 12'h509;
            14'd 3369: out = 12'h509;
            14'd 3370: out = 12'h509;
            14'd 3371: out = 12'h509;
            14'd 3372: out = 12'h509;
            14'd 3373: out = 12'h509;
            14'd 3374: out = 12'h50A;
            14'd 3375: out = 12'h50A;
            14'd 3376: out = 12'h50A;
            14'd 3377: out = 12'h50A;
            14'd 3378: out = 12'h50A;
            14'd 3379: out = 12'h50A;
            14'd 3380: out = 12'h50A;
            14'd 3381: out = 12'h50A;
            14'd 3382: out = 12'h50A;
            14'd 3383: out = 12'h50A;
            14'd 3384: out = 12'h50B;
            14'd 3385: out = 12'h50B;
            14'd 3386: out = 12'h50B;
            14'd 3387: out = 12'h50B;
            14'd 3388: out = 12'h50B;
            14'd 3389: out = 12'h50B;
            14'd 3390: out = 12'h50B;
            14'd 3391: out = 12'h50B;
            14'd 3392: out = 12'h50B;
            14'd 3393: out = 12'h50B;
            14'd 3394: out = 12'h50C;
            14'd 3395: out = 12'h50C;
            14'd 3396: out = 12'h50C;
            14'd 3397: out = 12'h50C;
            14'd 3398: out = 12'h50C;
            14'd 3399: out = 12'h50C;
            14'd 3400: out = 12'h50C;
            14'd 3401: out = 12'h50C;
            14'd 3402: out = 12'h50C;
            14'd 3403: out = 12'h50C;
            14'd 3404: out = 12'h50D;
            14'd 3405: out = 12'h50D;
            14'd 3406: out = 12'h50D;
            14'd 3407: out = 12'h50D;
            14'd 3408: out = 12'h50D;
            14'd 3409: out = 12'h50D;
            14'd 3410: out = 12'h50D;
            14'd 3411: out = 12'h50D;
            14'd 3412: out = 12'h50D;
            14'd 3413: out = 12'h50D;
            14'd 3414: out = 12'h50E;
            14'd 3415: out = 12'h50E;
            14'd 3416: out = 12'h50E;
            14'd 3417: out = 12'h50E;
            14'd 3418: out = 12'h50E;
            14'd 3419: out = 12'h50E;
            14'd 3420: out = 12'h50E;
            14'd 3421: out = 12'h50E;
            14'd 3422: out = 12'h50E;
            14'd 3423: out = 12'h50E;
            14'd 3424: out = 12'h50F;
            14'd 3425: out = 12'h50F;
            14'd 3426: out = 12'h50F;
            14'd 3427: out = 12'h50F;
            14'd 3428: out = 12'h50F;
            14'd 3429: out = 12'h50F;
            14'd 3430: out = 12'h50F;
            14'd 3431: out = 12'h50F;
            14'd 3432: out = 12'h50F;
            14'd 3433: out = 12'h50F;
            14'd 3434: out = 12'h510;
            14'd 3435: out = 12'h510;
            14'd 3436: out = 12'h510;
            14'd 3437: out = 12'h510;
            14'd 3438: out = 12'h510;
            14'd 3439: out = 12'h510;
            14'd 3440: out = 12'h510;
            14'd 3441: out = 12'h510;
            14'd 3442: out = 12'h510;
            14'd 3443: out = 12'h510;
            14'd 3444: out = 12'h511;
            14'd 3445: out = 12'h511;
            14'd 3446: out = 12'h511;
            14'd 3447: out = 12'h511;
            14'd 3448: out = 12'h511;
            14'd 3449: out = 12'h511;
            14'd 3450: out = 12'h511;
            14'd 3451: out = 12'h511;
            14'd 3452: out = 12'h511;
            14'd 3453: out = 12'h511;
            14'd 3454: out = 12'h512;
            14'd 3455: out = 12'h512;
            14'd 3456: out = 12'h512;
            14'd 3457: out = 12'h512;
            14'd 3458: out = 12'h512;
            14'd 3459: out = 12'h512;
            14'd 3460: out = 12'h512;
            14'd 3461: out = 12'h512;
            14'd 3462: out = 12'h512;
            14'd 3463: out = 12'h512;
            14'd 3464: out = 12'h513;
            14'd 3465: out = 12'h513;
            14'd 3466: out = 12'h513;
            14'd 3467: out = 12'h513;
            14'd 3468: out = 12'h513;
            14'd 3469: out = 12'h513;
            14'd 3470: out = 12'h513;
            14'd 3471: out = 12'h513;
            14'd 3472: out = 12'h513;
            14'd 3473: out = 12'h513;
            14'd 3474: out = 12'h514;
            14'd 3475: out = 12'h514;
            14'd 3476: out = 12'h514;
            14'd 3477: out = 12'h514;
            14'd 3478: out = 12'h514;
            14'd 3479: out = 12'h514;
            14'd 3480: out = 12'h514;
            14'd 3481: out = 12'h514;
            14'd 3482: out = 12'h514;
            14'd 3483: out = 12'h514;
            14'd 3484: out = 12'h515;
            14'd 3485: out = 12'h515;
            14'd 3486: out = 12'h515;
            14'd 3487: out = 12'h515;
            14'd 3488: out = 12'h515;
            14'd 3489: out = 12'h515;
            14'd 3490: out = 12'h515;
            14'd 3491: out = 12'h515;
            14'd 3492: out = 12'h515;
            14'd 3493: out = 12'h515;
            14'd 3494: out = 12'h516;
            14'd 3495: out = 12'h516;
            14'd 3496: out = 12'h516;
            14'd 3497: out = 12'h516;
            14'd 3498: out = 12'h516;
            14'd 3499: out = 12'h516;
            14'd 3500: out = 12'h516;
            14'd 3501: out = 12'h516;
            14'd 3502: out = 12'h516;
            14'd 3503: out = 12'h516;
            14'd 3504: out = 12'h517;
            14'd 3505: out = 12'h517;
            14'd 3506: out = 12'h517;
            14'd 3507: out = 12'h517;
            14'd 3508: out = 12'h517;
            14'd 3509: out = 12'h517;
            14'd 3510: out = 12'h517;
            14'd 3511: out = 12'h517;
            14'd 3512: out = 12'h517;
            14'd 3513: out = 12'h517;
            14'd 3514: out = 12'h518;
            14'd 3515: out = 12'h518;
            14'd 3516: out = 12'h518;
            14'd 3517: out = 12'h518;
            14'd 3518: out = 12'h518;
            14'd 3519: out = 12'h518;
            14'd 3520: out = 12'h518;
            14'd 3521: out = 12'h518;
            14'd 3522: out = 12'h518;
            14'd 3523: out = 12'h519;
            14'd 3524: out = 12'h519;
            14'd 3525: out = 12'h519;
            14'd 3526: out = 12'h519;
            14'd 3527: out = 12'h519;
            14'd 3528: out = 12'h519;
            14'd 3529: out = 12'h519;
            14'd 3530: out = 12'h519;
            14'd 3531: out = 12'h519;
            14'd 3532: out = 12'h519;
            14'd 3533: out = 12'h51A;
            14'd 3534: out = 12'h51A;
            14'd 3535: out = 12'h51A;
            14'd 3536: out = 12'h51A;
            14'd 3537: out = 12'h51A;
            14'd 3538: out = 12'h51A;
            14'd 3539: out = 12'h51A;
            14'd 3540: out = 12'h51A;
            14'd 3541: out = 12'h51A;
            14'd 3542: out = 12'h51A;
            14'd 3543: out = 12'h51B;
            14'd 3544: out = 12'h51B;
            14'd 3545: out = 12'h51B;
            14'd 3546: out = 12'h51B;
            14'd 3547: out = 12'h51B;
            14'd 3548: out = 12'h51B;
            14'd 3549: out = 12'h51B;
            14'd 3550: out = 12'h51B;
            14'd 3551: out = 12'h51B;
            14'd 3552: out = 12'h51B;
            14'd 3553: out = 12'h51C;
            14'd 3554: out = 12'h51C;
            14'd 3555: out = 12'h51C;
            14'd 3556: out = 12'h51C;
            14'd 3557: out = 12'h51C;
            14'd 3558: out = 12'h51C;
            14'd 3559: out = 12'h51C;
            14'd 3560: out = 12'h51C;
            14'd 3561: out = 12'h51C;
            14'd 3562: out = 12'h51C;
            14'd 3563: out = 12'h51D;
            14'd 3564: out = 12'h51D;
            14'd 3565: out = 12'h51D;
            14'd 3566: out = 12'h51D;
            14'd 3567: out = 12'h51D;
            14'd 3568: out = 12'h51D;
            14'd 3569: out = 12'h51D;
            14'd 3570: out = 12'h51D;
            14'd 3571: out = 12'h51D;
            14'd 3572: out = 12'h51D;
            14'd 3573: out = 12'h51E;
            14'd 3574: out = 12'h51E;
            14'd 3575: out = 12'h51E;
            14'd 3576: out = 12'h51E;
            14'd 3577: out = 12'h51E;
            14'd 3578: out = 12'h51E;
            14'd 3579: out = 12'h51E;
            14'd 3580: out = 12'h51E;
            14'd 3581: out = 12'h51E;
            14'd 3582: out = 12'h51F;
            14'd 3583: out = 12'h51F;
            14'd 3584: out = 12'h51F;
            14'd 3585: out = 12'h51F;
            14'd 3586: out = 12'h51F;
            14'd 3587: out = 12'h51F;
            14'd 3588: out = 12'h51F;
            14'd 3589: out = 12'h51F;
            14'd 3590: out = 12'h51F;
            14'd 3591: out = 12'h51F;
            14'd 3592: out = 12'h520;
            14'd 3593: out = 12'h520;
            14'd 3594: out = 12'h520;
            14'd 3595: out = 12'h520;
            14'd 3596: out = 12'h520;
            14'd 3597: out = 12'h520;
            14'd 3598: out = 12'h520;
            14'd 3599: out = 12'h520;
            14'd 3600: out = 12'h520;
            14'd 3601: out = 12'h520;
            14'd 3602: out = 12'h521;
            14'd 3603: out = 12'h521;
            14'd 3604: out = 12'h521;
            14'd 3605: out = 12'h521;
            14'd 3606: out = 12'h521;
            14'd 3607: out = 12'h521;
            14'd 3608: out = 12'h521;
            14'd 3609: out = 12'h521;
            14'd 3610: out = 12'h521;
            14'd 3611: out = 12'h521;
            14'd 3612: out = 12'h522;
            14'd 3613: out = 12'h522;
            14'd 3614: out = 12'h522;
            14'd 3615: out = 12'h522;
            14'd 3616: out = 12'h522;
            14'd 3617: out = 12'h522;
            14'd 3618: out = 12'h522;
            14'd 3619: out = 12'h522;
            14'd 3620: out = 12'h522;
            14'd 3621: out = 12'h523;
            14'd 3622: out = 12'h523;
            14'd 3623: out = 12'h523;
            14'd 3624: out = 12'h523;
            14'd 3625: out = 12'h523;
            14'd 3626: out = 12'h523;
            14'd 3627: out = 12'h523;
            14'd 3628: out = 12'h523;
            14'd 3629: out = 12'h523;
            14'd 3630: out = 12'h523;
            14'd 3631: out = 12'h524;
            14'd 3632: out = 12'h524;
            14'd 3633: out = 12'h524;
            14'd 3634: out = 12'h524;
            14'd 3635: out = 12'h524;
            14'd 3636: out = 12'h524;
            14'd 3637: out = 12'h524;
            14'd 3638: out = 12'h524;
            14'd 3639: out = 12'h524;
            14'd 3640: out = 12'h524;
            14'd 3641: out = 12'h525;
            14'd 3642: out = 12'h525;
            14'd 3643: out = 12'h525;
            14'd 3644: out = 12'h525;
            14'd 3645: out = 12'h525;
            14'd 3646: out = 12'h525;
            14'd 3647: out = 12'h525;
            14'd 3648: out = 12'h525;
            14'd 3649: out = 12'h525;
            14'd 3650: out = 12'h526;
            14'd 3651: out = 12'h526;
            14'd 3652: out = 12'h526;
            14'd 3653: out = 12'h526;
            14'd 3654: out = 12'h526;
            14'd 3655: out = 12'h526;
            14'd 3656: out = 12'h526;
            14'd 3657: out = 12'h526;
            14'd 3658: out = 12'h526;
            14'd 3659: out = 12'h526;
            14'd 3660: out = 12'h527;
            14'd 3661: out = 12'h527;
            14'd 3662: out = 12'h527;
            14'd 3663: out = 12'h527;
            14'd 3664: out = 12'h527;
            14'd 3665: out = 12'h527;
            14'd 3666: out = 12'h527;
            14'd 3667: out = 12'h527;
            14'd 3668: out = 12'h527;
            14'd 3669: out = 12'h527;
            14'd 3670: out = 12'h528;
            14'd 3671: out = 12'h528;
            14'd 3672: out = 12'h528;
            14'd 3673: out = 12'h528;
            14'd 3674: out = 12'h528;
            14'd 3675: out = 12'h528;
            14'd 3676: out = 12'h528;
            14'd 3677: out = 12'h528;
            14'd 3678: out = 12'h528;
            14'd 3679: out = 12'h529;
            14'd 3680: out = 12'h529;
            14'd 3681: out = 12'h529;
            14'd 3682: out = 12'h529;
            14'd 3683: out = 12'h529;
            14'd 3684: out = 12'h529;
            14'd 3685: out = 12'h529;
            14'd 3686: out = 12'h529;
            14'd 3687: out = 12'h529;
            14'd 3688: out = 12'h529;
            14'd 3689: out = 12'h52A;
            14'd 3690: out = 12'h52A;
            14'd 3691: out = 12'h52A;
            14'd 3692: out = 12'h52A;
            14'd 3693: out = 12'h52A;
            14'd 3694: out = 12'h52A;
            14'd 3695: out = 12'h52A;
            14'd 3696: out = 12'h52A;
            14'd 3697: out = 12'h52A;
            14'd 3698: out = 12'h52A;
            14'd 3699: out = 12'h52B;
            14'd 3700: out = 12'h52B;
            14'd 3701: out = 12'h52B;
            14'd 3702: out = 12'h52B;
            14'd 3703: out = 12'h52B;
            14'd 3704: out = 12'h52B;
            14'd 3705: out = 12'h52B;
            14'd 3706: out = 12'h52B;
            14'd 3707: out = 12'h52B;
            14'd 3708: out = 12'h52C;
            14'd 3709: out = 12'h52C;
            14'd 3710: out = 12'h52C;
            14'd 3711: out = 12'h52C;
            14'd 3712: out = 12'h52C;
            14'd 3713: out = 12'h52C;
            14'd 3714: out = 12'h52C;
            14'd 3715: out = 12'h52C;
            14'd 3716: out = 12'h52C;
            14'd 3717: out = 12'h52C;
            14'd 3718: out = 12'h52D;
            14'd 3719: out = 12'h52D;
            14'd 3720: out = 12'h52D;
            14'd 3721: out = 12'h52D;
            14'd 3722: out = 12'h52D;
            14'd 3723: out = 12'h52D;
            14'd 3724: out = 12'h52D;
            14'd 3725: out = 12'h52D;
            14'd 3726: out = 12'h52D;
            14'd 3727: out = 12'h52E;
            14'd 3728: out = 12'h52E;
            14'd 3729: out = 12'h52E;
            14'd 3730: out = 12'h52E;
            14'd 3731: out = 12'h52E;
            14'd 3732: out = 12'h52E;
            14'd 3733: out = 12'h52E;
            14'd 3734: out = 12'h52E;
            14'd 3735: out = 12'h52E;
            14'd 3736: out = 12'h52E;
            14'd 3737: out = 12'h52F;
            14'd 3738: out = 12'h52F;
            14'd 3739: out = 12'h52F;
            14'd 3740: out = 12'h52F;
            14'd 3741: out = 12'h52F;
            14'd 3742: out = 12'h52F;
            14'd 3743: out = 12'h52F;
            14'd 3744: out = 12'h52F;
            14'd 3745: out = 12'h52F;
            14'd 3746: out = 12'h530;
            14'd 3747: out = 12'h530;
            14'd 3748: out = 12'h530;
            14'd 3749: out = 12'h530;
            14'd 3750: out = 12'h530;
            14'd 3751: out = 12'h530;
            14'd 3752: out = 12'h530;
            14'd 3753: out = 12'h530;
            14'd 3754: out = 12'h530;
            14'd 3755: out = 12'h530;
            14'd 3756: out = 12'h531;
            14'd 3757: out = 12'h531;
            14'd 3758: out = 12'h531;
            14'd 3759: out = 12'h531;
            14'd 3760: out = 12'h531;
            14'd 3761: out = 12'h531;
            14'd 3762: out = 12'h531;
            14'd 3763: out = 12'h531;
            14'd 3764: out = 12'h531;
            14'd 3765: out = 12'h532;
            14'd 3766: out = 12'h532;
            14'd 3767: out = 12'h532;
            14'd 3768: out = 12'h532;
            14'd 3769: out = 12'h532;
            14'd 3770: out = 12'h532;
            14'd 3771: out = 12'h532;
            14'd 3772: out = 12'h532;
            14'd 3773: out = 12'h532;
            14'd 3774: out = 12'h532;
            14'd 3775: out = 12'h533;
            14'd 3776: out = 12'h533;
            14'd 3777: out = 12'h533;
            14'd 3778: out = 12'h533;
            14'd 3779: out = 12'h533;
            14'd 3780: out = 12'h533;
            14'd 3781: out = 12'h533;
            14'd 3782: out = 12'h533;
            14'd 3783: out = 12'h533;
            14'd 3784: out = 12'h534;
            14'd 3785: out = 12'h534;
            14'd 3786: out = 12'h534;
            14'd 3787: out = 12'h534;
            14'd 3788: out = 12'h534;
            14'd 3789: out = 12'h534;
            14'd 3790: out = 12'h534;
            14'd 3791: out = 12'h534;
            14'd 3792: out = 12'h534;
            14'd 3793: out = 12'h534;
            14'd 3794: out = 12'h535;
            14'd 3795: out = 12'h535;
            14'd 3796: out = 12'h535;
            14'd 3797: out = 12'h535;
            14'd 3798: out = 12'h535;
            14'd 3799: out = 12'h535;
            14'd 3800: out = 12'h535;
            14'd 3801: out = 12'h535;
            14'd 3802: out = 12'h535;
            14'd 3803: out = 12'h536;
            14'd 3804: out = 12'h536;
            14'd 3805: out = 12'h536;
            14'd 3806: out = 12'h536;
            14'd 3807: out = 12'h536;
            14'd 3808: out = 12'h536;
            14'd 3809: out = 12'h536;
            14'd 3810: out = 12'h536;
            14'd 3811: out = 12'h536;
            14'd 3812: out = 12'h536;
            14'd 3813: out = 12'h537;
            14'd 3814: out = 12'h537;
            14'd 3815: out = 12'h537;
            14'd 3816: out = 12'h537;
            14'd 3817: out = 12'h537;
            14'd 3818: out = 12'h537;
            14'd 3819: out = 12'h537;
            14'd 3820: out = 12'h537;
            14'd 3821: out = 12'h537;
            14'd 3822: out = 12'h538;
            14'd 3823: out = 12'h538;
            14'd 3824: out = 12'h538;
            14'd 3825: out = 12'h538;
            14'd 3826: out = 12'h538;
            14'd 3827: out = 12'h538;
            14'd 3828: out = 12'h538;
            14'd 3829: out = 12'h538;
            14'd 3830: out = 12'h538;
            14'd 3831: out = 12'h539;
            14'd 3832: out = 12'h539;
            14'd 3833: out = 12'h539;
            14'd 3834: out = 12'h539;
            14'd 3835: out = 12'h539;
            14'd 3836: out = 12'h539;
            14'd 3837: out = 12'h539;
            14'd 3838: out = 12'h539;
            14'd 3839: out = 12'h539;
            14'd 3840: out = 12'h539;
            14'd 3841: out = 12'h53A;
            14'd 3842: out = 12'h53A;
            14'd 3843: out = 12'h53A;
            14'd 3844: out = 12'h53A;
            14'd 3845: out = 12'h53A;
            14'd 3846: out = 12'h53A;
            14'd 3847: out = 12'h53A;
            14'd 3848: out = 12'h53A;
            14'd 3849: out = 12'h53A;
            14'd 3850: out = 12'h53B;
            14'd 3851: out = 12'h53B;
            14'd 3852: out = 12'h53B;
            14'd 3853: out = 12'h53B;
            14'd 3854: out = 12'h53B;
            14'd 3855: out = 12'h53B;
            14'd 3856: out = 12'h53B;
            14'd 3857: out = 12'h53B;
            14'd 3858: out = 12'h53B;
            14'd 3859: out = 12'h53B;
            14'd 3860: out = 12'h53C;
            14'd 3861: out = 12'h53C;
            14'd 3862: out = 12'h53C;
            14'd 3863: out = 12'h53C;
            14'd 3864: out = 12'h53C;
            14'd 3865: out = 12'h53C;
            14'd 3866: out = 12'h53C;
            14'd 3867: out = 12'h53C;
            14'd 3868: out = 12'h53C;
            14'd 3869: out = 12'h53D;
            14'd 3870: out = 12'h53D;
            14'd 3871: out = 12'h53D;
            14'd 3872: out = 12'h53D;
            14'd 3873: out = 12'h53D;
            14'd 3874: out = 12'h53D;
            14'd 3875: out = 12'h53D;
            14'd 3876: out = 12'h53D;
            14'd 3877: out = 12'h53D;
            14'd 3878: out = 12'h53E;
            14'd 3879: out = 12'h53E;
            14'd 3880: out = 12'h53E;
            14'd 3881: out = 12'h53E;
            14'd 3882: out = 12'h53E;
            14'd 3883: out = 12'h53E;
            14'd 3884: out = 12'h53E;
            14'd 3885: out = 12'h53E;
            14'd 3886: out = 12'h53E;
            14'd 3887: out = 12'h53E;
            14'd 3888: out = 12'h53F;
            14'd 3889: out = 12'h53F;
            14'd 3890: out = 12'h53F;
            14'd 3891: out = 12'h53F;
            14'd 3892: out = 12'h53F;
            14'd 3893: out = 12'h53F;
            14'd 3894: out = 12'h53F;
            14'd 3895: out = 12'h53F;
            14'd 3896: out = 12'h53F;
            14'd 3897: out = 12'h540;
            14'd 3898: out = 12'h540;
            14'd 3899: out = 12'h540;
            14'd 3900: out = 12'h540;
            14'd 3901: out = 12'h540;
            14'd 3902: out = 12'h540;
            14'd 3903: out = 12'h540;
            14'd 3904: out = 12'h540;
            14'd 3905: out = 12'h540;
            14'd 3906: out = 12'h541;
            14'd 3907: out = 12'h541;
            14'd 3908: out = 12'h541;
            14'd 3909: out = 12'h541;
            14'd 3910: out = 12'h541;
            14'd 3911: out = 12'h541;
            14'd 3912: out = 12'h541;
            14'd 3913: out = 12'h541;
            14'd 3914: out = 12'h541;
            14'd 3915: out = 12'h542;
            14'd 3916: out = 12'h542;
            14'd 3917: out = 12'h542;
            14'd 3918: out = 12'h542;
            14'd 3919: out = 12'h542;
            14'd 3920: out = 12'h542;
            14'd 3921: out = 12'h542;
            14'd 3922: out = 12'h542;
            14'd 3923: out = 12'h542;
            14'd 3924: out = 12'h542;
            14'd 3925: out = 12'h543;
            14'd 3926: out = 12'h543;
            14'd 3927: out = 12'h543;
            14'd 3928: out = 12'h543;
            14'd 3929: out = 12'h543;
            14'd 3930: out = 12'h543;
            14'd 3931: out = 12'h543;
            14'd 3932: out = 12'h543;
            14'd 3933: out = 12'h543;
            14'd 3934: out = 12'h544;
            14'd 3935: out = 12'h544;
            14'd 3936: out = 12'h544;
            14'd 3937: out = 12'h544;
            14'd 3938: out = 12'h544;
            14'd 3939: out = 12'h544;
            14'd 3940: out = 12'h544;
            14'd 3941: out = 12'h544;
            14'd 3942: out = 12'h544;
            14'd 3943: out = 12'h545;
            14'd 3944: out = 12'h545;
            14'd 3945: out = 12'h545;
            14'd 3946: out = 12'h545;
            14'd 3947: out = 12'h545;
            14'd 3948: out = 12'h545;
            14'd 3949: out = 12'h545;
            14'd 3950: out = 12'h545;
            14'd 3951: out = 12'h545;
            14'd 3952: out = 12'h546;
            14'd 3953: out = 12'h546;
            14'd 3954: out = 12'h546;
            14'd 3955: out = 12'h546;
            14'd 3956: out = 12'h546;
            14'd 3957: out = 12'h546;
            14'd 3958: out = 12'h546;
            14'd 3959: out = 12'h546;
            14'd 3960: out = 12'h546;
            14'd 3961: out = 12'h546;
            14'd 3962: out = 12'h547;
            14'd 3963: out = 12'h547;
            14'd 3964: out = 12'h547;
            14'd 3965: out = 12'h547;
            14'd 3966: out = 12'h547;
            14'd 3967: out = 12'h547;
            14'd 3968: out = 12'h547;
            14'd 3969: out = 12'h547;
            14'd 3970: out = 12'h547;
            14'd 3971: out = 12'h548;
            14'd 3972: out = 12'h548;
            14'd 3973: out = 12'h548;
            14'd 3974: out = 12'h548;
            14'd 3975: out = 12'h548;
            14'd 3976: out = 12'h548;
            14'd 3977: out = 12'h548;
            14'd 3978: out = 12'h548;
            14'd 3979: out = 12'h548;
            14'd 3980: out = 12'h549;
            14'd 3981: out = 12'h549;
            14'd 3982: out = 12'h549;
            14'd 3983: out = 12'h549;
            14'd 3984: out = 12'h549;
            14'd 3985: out = 12'h549;
            14'd 3986: out = 12'h549;
            14'd 3987: out = 12'h549;
            14'd 3988: out = 12'h549;
            14'd 3989: out = 12'h54A;
            14'd 3990: out = 12'h54A;
            14'd 3991: out = 12'h54A;
            14'd 3992: out = 12'h54A;
            14'd 3993: out = 12'h54A;
            14'd 3994: out = 12'h54A;
            14'd 3995: out = 12'h54A;
            14'd 3996: out = 12'h54A;
            14'd 3997: out = 12'h54A;
            14'd 3998: out = 12'h54B;
            14'd 3999: out = 12'h54B;
            14'd 4000: out = 12'h54B;
            14'd 4001: out = 12'h54B;
            14'd 4002: out = 12'h54B;
            14'd 4003: out = 12'h54B;
            14'd 4004: out = 12'h54B;
            14'd 4005: out = 12'h54B;
            14'd 4006: out = 12'h54B;
            14'd 4007: out = 12'h54C;
            14'd 4008: out = 12'h54C;
            14'd 4009: out = 12'h54C;
            14'd 4010: out = 12'h54C;
            14'd 4011: out = 12'h54C;
            14'd 4012: out = 12'h54C;
            14'd 4013: out = 12'h54C;
            14'd 4014: out = 12'h54C;
            14'd 4015: out = 12'h54C;
            14'd 4016: out = 12'h54D;
            14'd 4017: out = 12'h54D;
            14'd 4018: out = 12'h54D;
            14'd 4019: out = 12'h54D;
            14'd 4020: out = 12'h54D;
            14'd 4021: out = 12'h54D;
            14'd 4022: out = 12'h54D;
            14'd 4023: out = 12'h54D;
            14'd 4024: out = 12'h54D;
            14'd 4025: out = 12'h54D;
            14'd 4026: out = 12'h54E;
            14'd 4027: out = 12'h54E;
            14'd 4028: out = 12'h54E;
            14'd 4029: out = 12'h54E;
            14'd 4030: out = 12'h54E;
            14'd 4031: out = 12'h54E;
            14'd 4032: out = 12'h54E;
            14'd 4033: out = 12'h54E;
            14'd 4034: out = 12'h54E;
            14'd 4035: out = 12'h54F;
            14'd 4036: out = 12'h54F;
            14'd 4037: out = 12'h54F;
            14'd 4038: out = 12'h54F;
            14'd 4039: out = 12'h54F;
            14'd 4040: out = 12'h54F;
            14'd 4041: out = 12'h54F;
            14'd 4042: out = 12'h54F;
            14'd 4043: out = 12'h54F;
            14'd 4044: out = 12'h550;
            14'd 4045: out = 12'h550;
            14'd 4046: out = 12'h550;
            14'd 4047: out = 12'h550;
            14'd 4048: out = 12'h550;
            14'd 4049: out = 12'h550;
            14'd 4050: out = 12'h550;
            14'd 4051: out = 12'h550;
            14'd 4052: out = 12'h550;
            14'd 4053: out = 12'h551;
            14'd 4054: out = 12'h551;
            14'd 4055: out = 12'h551;
            14'd 4056: out = 12'h551;
            14'd 4057: out = 12'h551;
            14'd 4058: out = 12'h551;
            14'd 4059: out = 12'h551;
            14'd 4060: out = 12'h551;
            14'd 4061: out = 12'h551;
            14'd 4062: out = 12'h552;
            14'd 4063: out = 12'h552;
            14'd 4064: out = 12'h552;
            14'd 4065: out = 12'h552;
            14'd 4066: out = 12'h552;
            14'd 4067: out = 12'h552;
            14'd 4068: out = 12'h552;
            14'd 4069: out = 12'h552;
            14'd 4070: out = 12'h552;
            14'd 4071: out = 12'h553;
            14'd 4072: out = 12'h553;
            14'd 4073: out = 12'h553;
            14'd 4074: out = 12'h553;
            14'd 4075: out = 12'h553;
            14'd 4076: out = 12'h553;
            14'd 4077: out = 12'h553;
            14'd 4078: out = 12'h553;
            14'd 4079: out = 12'h553;
            14'd 4080: out = 12'h554;
            14'd 4081: out = 12'h554;
            14'd 4082: out = 12'h554;
            14'd 4083: out = 12'h554;
            14'd 4084: out = 12'h554;
            14'd 4085: out = 12'h554;
            14'd 4086: out = 12'h554;
            14'd 4087: out = 12'h554;
            14'd 4088: out = 12'h554;
            14'd 4089: out = 12'h555;
            14'd 4090: out = 12'h555;
            14'd 4091: out = 12'h555;
            14'd 4092: out = 12'h555;
            14'd 4093: out = 12'h555;
            14'd 4094: out = 12'h555;
            14'd 4095: out = 12'h555;
            14'd 4096: out = 12'h555;
            14'd 4097: out = 12'h555;
            14'd 4098: out = 12'h556;
            14'd 4099: out = 12'h556;
            14'd 4100: out = 12'h556;
            14'd 4101: out = 12'h556;
            14'd 4102: out = 12'h556;
            14'd 4103: out = 12'h556;
            14'd 4104: out = 12'h556;
            14'd 4105: out = 12'h556;
            14'd 4106: out = 12'h556;
            14'd 4107: out = 12'h557;
            14'd 4108: out = 12'h557;
            14'd 4109: out = 12'h557;
            14'd 4110: out = 12'h557;
            14'd 4111: out = 12'h557;
            14'd 4112: out = 12'h557;
            14'd 4113: out = 12'h557;
            14'd 4114: out = 12'h557;
            14'd 4115: out = 12'h557;
            14'd 4116: out = 12'h558;
            14'd 4117: out = 12'h558;
            14'd 4118: out = 12'h558;
            14'd 4119: out = 12'h558;
            14'd 4120: out = 12'h558;
            14'd 4121: out = 12'h558;
            14'd 4122: out = 12'h558;
            14'd 4123: out = 12'h558;
            14'd 4124: out = 12'h558;
            14'd 4125: out = 12'h559;
            14'd 4126: out = 12'h559;
            14'd 4127: out = 12'h559;
            14'd 4128: out = 12'h559;
            14'd 4129: out = 12'h559;
            14'd 4130: out = 12'h559;
            14'd 4131: out = 12'h559;
            14'd 4132: out = 12'h559;
            14'd 4133: out = 12'h559;
            14'd 4134: out = 12'h55A;
            14'd 4135: out = 12'h55A;
            14'd 4136: out = 12'h55A;
            14'd 4137: out = 12'h55A;
            14'd 4138: out = 12'h55A;
            14'd 4139: out = 12'h55A;
            14'd 4140: out = 12'h55A;
            14'd 4141: out = 12'h55A;
            14'd 4142: out = 12'h55A;
            14'd 4143: out = 12'h55B;
            14'd 4144: out = 12'h55B;
            14'd 4145: out = 12'h55B;
            14'd 4146: out = 12'h55B;
            14'd 4147: out = 12'h55B;
            14'd 4148: out = 12'h55B;
            14'd 4149: out = 12'h55B;
            14'd 4150: out = 12'h55B;
            14'd 4151: out = 12'h55B;
            14'd 4152: out = 12'h55C;
            14'd 4153: out = 12'h55C;
            14'd 4154: out = 12'h55C;
            14'd 4155: out = 12'h55C;
            14'd 4156: out = 12'h55C;
            14'd 4157: out = 12'h55C;
            14'd 4158: out = 12'h55C;
            14'd 4159: out = 12'h55C;
            14'd 4160: out = 12'h55C;
            14'd 4161: out = 12'h55D;
            14'd 4162: out = 12'h55D;
            14'd 4163: out = 12'h55D;
            14'd 4164: out = 12'h55D;
            14'd 4165: out = 12'h55D;
            14'd 4166: out = 12'h55D;
            14'd 4167: out = 12'h55D;
            14'd 4168: out = 12'h55D;
            14'd 4169: out = 12'h55D;
            14'd 4170: out = 12'h55E;
            14'd 4171: out = 12'h55E;
            14'd 4172: out = 12'h55E;
            14'd 4173: out = 12'h55E;
            14'd 4174: out = 12'h55E;
            14'd 4175: out = 12'h55E;
            14'd 4176: out = 12'h55E;
            14'd 4177: out = 12'h55E;
            14'd 4178: out = 12'h55F;
            14'd 4179: out = 12'h55F;
            14'd 4180: out = 12'h55F;
            14'd 4181: out = 12'h55F;
            14'd 4182: out = 12'h55F;
            14'd 4183: out = 12'h55F;
            14'd 4184: out = 12'h55F;
            14'd 4185: out = 12'h55F;
            14'd 4186: out = 12'h55F;
            14'd 4187: out = 12'h560;
            14'd 4188: out = 12'h560;
            14'd 4189: out = 12'h560;
            14'd 4190: out = 12'h560;
            14'd 4191: out = 12'h560;
            14'd 4192: out = 12'h560;
            14'd 4193: out = 12'h560;
            14'd 4194: out = 12'h560;
            14'd 4195: out = 12'h560;
            14'd 4196: out = 12'h561;
            14'd 4197: out = 12'h561;
            14'd 4198: out = 12'h561;
            14'd 4199: out = 12'h561;
            14'd 4200: out = 12'h561;
            14'd 4201: out = 12'h561;
            14'd 4202: out = 12'h561;
            14'd 4203: out = 12'h561;
            14'd 4204: out = 12'h561;
            14'd 4205: out = 12'h562;
            14'd 4206: out = 12'h562;
            14'd 4207: out = 12'h562;
            14'd 4208: out = 12'h562;
            14'd 4209: out = 12'h562;
            14'd 4210: out = 12'h562;
            14'd 4211: out = 12'h562;
            14'd 4212: out = 12'h562;
            14'd 4213: out = 12'h562;
            14'd 4214: out = 12'h563;
            14'd 4215: out = 12'h563;
            14'd 4216: out = 12'h563;
            14'd 4217: out = 12'h563;
            14'd 4218: out = 12'h563;
            14'd 4219: out = 12'h563;
            14'd 4220: out = 12'h563;
            14'd 4221: out = 12'h563;
            14'd 4222: out = 12'h563;
            14'd 4223: out = 12'h564;
            14'd 4224: out = 12'h564;
            14'd 4225: out = 12'h564;
            14'd 4226: out = 12'h564;
            14'd 4227: out = 12'h564;
            14'd 4228: out = 12'h564;
            14'd 4229: out = 12'h564;
            14'd 4230: out = 12'h564;
            14'd 4231: out = 12'h564;
            14'd 4232: out = 12'h565;
            14'd 4233: out = 12'h565;
            14'd 4234: out = 12'h565;
            14'd 4235: out = 12'h565;
            14'd 4236: out = 12'h565;
            14'd 4237: out = 12'h565;
            14'd 4238: out = 12'h565;
            14'd 4239: out = 12'h565;
            14'd 4240: out = 12'h566;
            14'd 4241: out = 12'h566;
            14'd 4242: out = 12'h566;
            14'd 4243: out = 12'h566;
            14'd 4244: out = 12'h566;
            14'd 4245: out = 12'h566;
            14'd 4246: out = 12'h566;
            14'd 4247: out = 12'h566;
            14'd 4248: out = 12'h566;
            14'd 4249: out = 12'h567;
            14'd 4250: out = 12'h567;
            14'd 4251: out = 12'h567;
            14'd 4252: out = 12'h567;
            14'd 4253: out = 12'h567;
            14'd 4254: out = 12'h567;
            14'd 4255: out = 12'h567;
            14'd 4256: out = 12'h567;
            14'd 4257: out = 12'h567;
            14'd 4258: out = 12'h568;
            14'd 4259: out = 12'h568;
            14'd 4260: out = 12'h568;
            14'd 4261: out = 12'h568;
            14'd 4262: out = 12'h568;
            14'd 4263: out = 12'h568;
            14'd 4264: out = 12'h568;
            14'd 4265: out = 12'h568;
            14'd 4266: out = 12'h568;
            14'd 4267: out = 12'h569;
            14'd 4268: out = 12'h569;
            14'd 4269: out = 12'h569;
            14'd 4270: out = 12'h569;
            14'd 4271: out = 12'h569;
            14'd 4272: out = 12'h569;
            14'd 4273: out = 12'h569;
            14'd 4274: out = 12'h569;
            14'd 4275: out = 12'h56A;
            14'd 4276: out = 12'h56A;
            14'd 4277: out = 12'h56A;
            14'd 4278: out = 12'h56A;
            14'd 4279: out = 12'h56A;
            14'd 4280: out = 12'h56A;
            14'd 4281: out = 12'h56A;
            14'd 4282: out = 12'h56A;
            14'd 4283: out = 12'h56A;
            14'd 4284: out = 12'h56B;
            14'd 4285: out = 12'h56B;
            14'd 4286: out = 12'h56B;
            14'd 4287: out = 12'h56B;
            14'd 4288: out = 12'h56B;
            14'd 4289: out = 12'h56B;
            14'd 4290: out = 12'h56B;
            14'd 4291: out = 12'h56B;
            14'd 4292: out = 12'h56B;
            14'd 4293: out = 12'h56C;
            14'd 4294: out = 12'h56C;
            14'd 4295: out = 12'h56C;
            14'd 4296: out = 12'h56C;
            14'd 4297: out = 12'h56C;
            14'd 4298: out = 12'h56C;
            14'd 4299: out = 12'h56C;
            14'd 4300: out = 12'h56C;
            14'd 4301: out = 12'h56C;
            14'd 4302: out = 12'h56D;
            14'd 4303: out = 12'h56D;
            14'd 4304: out = 12'h56D;
            14'd 4305: out = 12'h56D;
            14'd 4306: out = 12'h56D;
            14'd 4307: out = 12'h56D;
            14'd 4308: out = 12'h56D;
            14'd 4309: out = 12'h56D;
            14'd 4310: out = 12'h56E;
            14'd 4311: out = 12'h56E;
            14'd 4312: out = 12'h56E;
            14'd 4313: out = 12'h56E;
            14'd 4314: out = 12'h56E;
            14'd 4315: out = 12'h56E;
            14'd 4316: out = 12'h56E;
            14'd 4317: out = 12'h56E;
            14'd 4318: out = 12'h56E;
            14'd 4319: out = 12'h56F;
            14'd 4320: out = 12'h56F;
            14'd 4321: out = 12'h56F;
            14'd 4322: out = 12'h56F;
            14'd 4323: out = 12'h56F;
            14'd 4324: out = 12'h56F;
            14'd 4325: out = 12'h56F;
            14'd 4326: out = 12'h56F;
            14'd 4327: out = 12'h56F;
            14'd 4328: out = 12'h570;
            14'd 4329: out = 12'h570;
            14'd 4330: out = 12'h570;
            14'd 4331: out = 12'h570;
            14'd 4332: out = 12'h570;
            14'd 4333: out = 12'h570;
            14'd 4334: out = 12'h570;
            14'd 4335: out = 12'h570;
            14'd 4336: out = 12'h571;
            14'd 4337: out = 12'h571;
            14'd 4338: out = 12'h571;
            14'd 4339: out = 12'h571;
            14'd 4340: out = 12'h571;
            14'd 4341: out = 12'h571;
            14'd 4342: out = 12'h571;
            14'd 4343: out = 12'h571;
            14'd 4344: out = 12'h571;
            14'd 4345: out = 12'h572;
            14'd 4346: out = 12'h572;
            14'd 4347: out = 12'h572;
            14'd 4348: out = 12'h572;
            14'd 4349: out = 12'h572;
            14'd 4350: out = 12'h572;
            14'd 4351: out = 12'h572;
            14'd 4352: out = 12'h572;
            14'd 4353: out = 12'h572;
            14'd 4354: out = 12'h573;
            14'd 4355: out = 12'h573;
            14'd 4356: out = 12'h573;
            14'd 4357: out = 12'h573;
            14'd 4358: out = 12'h573;
            14'd 4359: out = 12'h573;
            14'd 4360: out = 12'h573;
            14'd 4361: out = 12'h573;
            14'd 4362: out = 12'h574;
            14'd 4363: out = 12'h574;
            14'd 4364: out = 12'h574;
            14'd 4365: out = 12'h574;
            14'd 4366: out = 12'h574;
            14'd 4367: out = 12'h574;
            14'd 4368: out = 12'h574;
            14'd 4369: out = 12'h574;
            14'd 4370: out = 12'h574;
            14'd 4371: out = 12'h575;
            14'd 4372: out = 12'h575;
            14'd 4373: out = 12'h575;
            14'd 4374: out = 12'h575;
            14'd 4375: out = 12'h575;
            14'd 4376: out = 12'h575;
            14'd 4377: out = 12'h575;
            14'd 4378: out = 12'h575;
            14'd 4379: out = 12'h576;
            14'd 4380: out = 12'h576;
            14'd 4381: out = 12'h576;
            14'd 4382: out = 12'h576;
            14'd 4383: out = 12'h576;
            14'd 4384: out = 12'h576;
            14'd 4385: out = 12'h576;
            14'd 4386: out = 12'h576;
            14'd 4387: out = 12'h576;
            14'd 4388: out = 12'h577;
            14'd 4389: out = 12'h577;
            14'd 4390: out = 12'h577;
            14'd 4391: out = 12'h577;
            14'd 4392: out = 12'h577;
            14'd 4393: out = 12'h577;
            14'd 4394: out = 12'h577;
            14'd 4395: out = 12'h577;
            14'd 4396: out = 12'h578;
            14'd 4397: out = 12'h578;
            14'd 4398: out = 12'h578;
            14'd 4399: out = 12'h578;
            14'd 4400: out = 12'h578;
            14'd 4401: out = 12'h578;
            14'd 4402: out = 12'h578;
            14'd 4403: out = 12'h578;
            14'd 4404: out = 12'h578;
            14'd 4405: out = 12'h579;
            14'd 4406: out = 12'h579;
            14'd 4407: out = 12'h579;
            14'd 4408: out = 12'h579;
            14'd 4409: out = 12'h579;
            14'd 4410: out = 12'h579;
            14'd 4411: out = 12'h579;
            14'd 4412: out = 12'h579;
            14'd 4413: out = 12'h579;
            14'd 4414: out = 12'h57A;
            14'd 4415: out = 12'h57A;
            14'd 4416: out = 12'h57A;
            14'd 4417: out = 12'h57A;
            14'd 4418: out = 12'h57A;
            14'd 4419: out = 12'h57A;
            14'd 4420: out = 12'h57A;
            14'd 4421: out = 12'h57A;
            14'd 4422: out = 12'h57B;
            14'd 4423: out = 12'h57B;
            14'd 4424: out = 12'h57B;
            14'd 4425: out = 12'h57B;
            14'd 4426: out = 12'h57B;
            14'd 4427: out = 12'h57B;
            14'd 4428: out = 12'h57B;
            14'd 4429: out = 12'h57B;
            14'd 4430: out = 12'h57B;
            14'd 4431: out = 12'h57C;
            14'd 4432: out = 12'h57C;
            14'd 4433: out = 12'h57C;
            14'd 4434: out = 12'h57C;
            14'd 4435: out = 12'h57C;
            14'd 4436: out = 12'h57C;
            14'd 4437: out = 12'h57C;
            14'd 4438: out = 12'h57C;
            14'd 4439: out = 12'h57D;
            14'd 4440: out = 12'h57D;
            14'd 4441: out = 12'h57D;
            14'd 4442: out = 12'h57D;
            14'd 4443: out = 12'h57D;
            14'd 4444: out = 12'h57D;
            14'd 4445: out = 12'h57D;
            14'd 4446: out = 12'h57D;
            14'd 4447: out = 12'h57D;
            14'd 4448: out = 12'h57E;
            14'd 4449: out = 12'h57E;
            14'd 4450: out = 12'h57E;
            14'd 4451: out = 12'h57E;
            14'd 4452: out = 12'h57E;
            14'd 4453: out = 12'h57E;
            14'd 4454: out = 12'h57E;
            14'd 4455: out = 12'h57E;
            14'd 4456: out = 12'h57F;
            14'd 4457: out = 12'h57F;
            14'd 4458: out = 12'h57F;
            14'd 4459: out = 12'h57F;
            14'd 4460: out = 12'h57F;
            14'd 4461: out = 12'h57F;
            14'd 4462: out = 12'h57F;
            14'd 4463: out = 12'h57F;
            14'd 4464: out = 12'h57F;
            14'd 4465: out = 12'h580;
            14'd 4466: out = 12'h580;
            14'd 4467: out = 12'h580;
            14'd 4468: out = 12'h580;
            14'd 4469: out = 12'h580;
            14'd 4470: out = 12'h580;
            14'd 4471: out = 12'h580;
            14'd 4472: out = 12'h580;
            14'd 4473: out = 12'h581;
            14'd 4474: out = 12'h581;
            14'd 4475: out = 12'h581;
            14'd 4476: out = 12'h581;
            14'd 4477: out = 12'h581;
            14'd 4478: out = 12'h581;
            14'd 4479: out = 12'h581;
            14'd 4480: out = 12'h581;
            14'd 4481: out = 12'h581;
            14'd 4482: out = 12'h582;
            14'd 4483: out = 12'h582;
            14'd 4484: out = 12'h582;
            14'd 4485: out = 12'h582;
            14'd 4486: out = 12'h582;
            14'd 4487: out = 12'h582;
            14'd 4488: out = 12'h582;
            14'd 4489: out = 12'h582;
            14'd 4490: out = 12'h583;
            14'd 4491: out = 12'h583;
            14'd 4492: out = 12'h583;
            14'd 4493: out = 12'h583;
            14'd 4494: out = 12'h583;
            14'd 4495: out = 12'h583;
            14'd 4496: out = 12'h583;
            14'd 4497: out = 12'h583;
            14'd 4498: out = 12'h584;
            14'd 4499: out = 12'h584;
            14'd 4500: out = 12'h584;
            14'd 4501: out = 12'h584;
            14'd 4502: out = 12'h584;
            14'd 4503: out = 12'h584;
            14'd 4504: out = 12'h584;
            14'd 4505: out = 12'h584;
            14'd 4506: out = 12'h584;
            14'd 4507: out = 12'h585;
            14'd 4508: out = 12'h585;
            14'd 4509: out = 12'h585;
            14'd 4510: out = 12'h585;
            14'd 4511: out = 12'h585;
            14'd 4512: out = 12'h585;
            14'd 4513: out = 12'h585;
            14'd 4514: out = 12'h585;
            14'd 4515: out = 12'h586;
            14'd 4516: out = 12'h586;
            14'd 4517: out = 12'h586;
            14'd 4518: out = 12'h586;
            14'd 4519: out = 12'h586;
            14'd 4520: out = 12'h586;
            14'd 4521: out = 12'h586;
            14'd 4522: out = 12'h586;
            14'd 4523: out = 12'h586;
            14'd 4524: out = 12'h587;
            14'd 4525: out = 12'h587;
            14'd 4526: out = 12'h587;
            14'd 4527: out = 12'h587;
            14'd 4528: out = 12'h587;
            14'd 4529: out = 12'h587;
            14'd 4530: out = 12'h587;
            14'd 4531: out = 12'h587;
            14'd 4532: out = 12'h588;
            14'd 4533: out = 12'h588;
            14'd 4534: out = 12'h588;
            14'd 4535: out = 12'h588;
            14'd 4536: out = 12'h588;
            14'd 4537: out = 12'h588;
            14'd 4538: out = 12'h588;
            14'd 4539: out = 12'h588;
            14'd 4540: out = 12'h589;
            14'd 4541: out = 12'h589;
            14'd 4542: out = 12'h589;
            14'd 4543: out = 12'h589;
            14'd 4544: out = 12'h589;
            14'd 4545: out = 12'h589;
            14'd 4546: out = 12'h589;
            14'd 4547: out = 12'h589;
            14'd 4548: out = 12'h589;
            14'd 4549: out = 12'h58A;
            14'd 4550: out = 12'h58A;
            14'd 4551: out = 12'h58A;
            14'd 4552: out = 12'h58A;
            14'd 4553: out = 12'h58A;
            14'd 4554: out = 12'h58A;
            14'd 4555: out = 12'h58A;
            14'd 4556: out = 12'h58A;
            14'd 4557: out = 12'h58B;
            14'd 4558: out = 12'h58B;
            14'd 4559: out = 12'h58B;
            14'd 4560: out = 12'h58B;
            14'd 4561: out = 12'h58B;
            14'd 4562: out = 12'h58B;
            14'd 4563: out = 12'h58B;
            14'd 4564: out = 12'h58B;
            14'd 4565: out = 12'h58C;
            14'd 4566: out = 12'h58C;
            14'd 4567: out = 12'h58C;
            14'd 4568: out = 12'h58C;
            14'd 4569: out = 12'h58C;
            14'd 4570: out = 12'h58C;
            14'd 4571: out = 12'h58C;
            14'd 4572: out = 12'h58C;
            14'd 4573: out = 12'h58C;
            14'd 4574: out = 12'h58D;
            14'd 4575: out = 12'h58D;
            14'd 4576: out = 12'h58D;
            14'd 4577: out = 12'h58D;
            14'd 4578: out = 12'h58D;
            14'd 4579: out = 12'h58D;
            14'd 4580: out = 12'h58D;
            14'd 4581: out = 12'h58D;
            14'd 4582: out = 12'h58E;
            14'd 4583: out = 12'h58E;
            14'd 4584: out = 12'h58E;
            14'd 4585: out = 12'h58E;
            14'd 4586: out = 12'h58E;
            14'd 4587: out = 12'h58E;
            14'd 4588: out = 12'h58E;
            14'd 4589: out = 12'h58E;
            14'd 4590: out = 12'h58F;
            14'd 4591: out = 12'h58F;
            14'd 4592: out = 12'h58F;
            14'd 4593: out = 12'h58F;
            14'd 4594: out = 12'h58F;
            14'd 4595: out = 12'h58F;
            14'd 4596: out = 12'h58F;
            14'd 4597: out = 12'h58F;
            14'd 4598: out = 12'h58F;
            14'd 4599: out = 12'h590;
            14'd 4600: out = 12'h590;
            14'd 4601: out = 12'h590;
            14'd 4602: out = 12'h590;
            14'd 4603: out = 12'h590;
            14'd 4604: out = 12'h590;
            14'd 4605: out = 12'h590;
            14'd 4606: out = 12'h590;
            14'd 4607: out = 12'h591;
            14'd 4608: out = 12'h591;
            14'd 4609: out = 12'h591;
            14'd 4610: out = 12'h591;
            14'd 4611: out = 12'h591;
            14'd 4612: out = 12'h591;
            14'd 4613: out = 12'h591;
            14'd 4614: out = 12'h591;
            14'd 4615: out = 12'h592;
            14'd 4616: out = 12'h592;
            14'd 4617: out = 12'h592;
            14'd 4618: out = 12'h592;
            14'd 4619: out = 12'h592;
            14'd 4620: out = 12'h592;
            14'd 4621: out = 12'h592;
            14'd 4622: out = 12'h592;
            14'd 4623: out = 12'h593;
            14'd 4624: out = 12'h593;
            14'd 4625: out = 12'h593;
            14'd 4626: out = 12'h593;
            14'd 4627: out = 12'h593;
            14'd 4628: out = 12'h593;
            14'd 4629: out = 12'h593;
            14'd 4630: out = 12'h593;
            14'd 4631: out = 12'h593;
            14'd 4632: out = 12'h594;
            14'd 4633: out = 12'h594;
            14'd 4634: out = 12'h594;
            14'd 4635: out = 12'h594;
            14'd 4636: out = 12'h594;
            14'd 4637: out = 12'h594;
            14'd 4638: out = 12'h594;
            14'd 4639: out = 12'h594;
            14'd 4640: out = 12'h595;
            14'd 4641: out = 12'h595;
            14'd 4642: out = 12'h595;
            14'd 4643: out = 12'h595;
            14'd 4644: out = 12'h595;
            14'd 4645: out = 12'h595;
            14'd 4646: out = 12'h595;
            14'd 4647: out = 12'h595;
            14'd 4648: out = 12'h596;
            14'd 4649: out = 12'h596;
            14'd 4650: out = 12'h596;
            14'd 4651: out = 12'h596;
            14'd 4652: out = 12'h596;
            14'd 4653: out = 12'h596;
            14'd 4654: out = 12'h596;
            14'd 4655: out = 12'h596;
            14'd 4656: out = 12'h597;
            14'd 4657: out = 12'h597;
            14'd 4658: out = 12'h597;
            14'd 4659: out = 12'h597;
            14'd 4660: out = 12'h597;
            14'd 4661: out = 12'h597;
            14'd 4662: out = 12'h597;
            14'd 4663: out = 12'h597;
            14'd 4664: out = 12'h598;
            14'd 4665: out = 12'h598;
            14'd 4666: out = 12'h598;
            14'd 4667: out = 12'h598;
            14'd 4668: out = 12'h598;
            14'd 4669: out = 12'h598;
            14'd 4670: out = 12'h598;
            14'd 4671: out = 12'h598;
            14'd 4672: out = 12'h598;
            14'd 4673: out = 12'h599;
            14'd 4674: out = 12'h599;
            14'd 4675: out = 12'h599;
            14'd 4676: out = 12'h599;
            14'd 4677: out = 12'h599;
            14'd 4678: out = 12'h599;
            14'd 4679: out = 12'h599;
            14'd 4680: out = 12'h599;
            14'd 4681: out = 12'h59A;
            14'd 4682: out = 12'h59A;
            14'd 4683: out = 12'h59A;
            14'd 4684: out = 12'h59A;
            14'd 4685: out = 12'h59A;
            14'd 4686: out = 12'h59A;
            14'd 4687: out = 12'h59A;
            14'd 4688: out = 12'h59A;
            14'd 4689: out = 12'h59B;
            14'd 4690: out = 12'h59B;
            14'd 4691: out = 12'h59B;
            14'd 4692: out = 12'h59B;
            14'd 4693: out = 12'h59B;
            14'd 4694: out = 12'h59B;
            14'd 4695: out = 12'h59B;
            14'd 4696: out = 12'h59B;
            14'd 4697: out = 12'h59C;
            14'd 4698: out = 12'h59C;
            14'd 4699: out = 12'h59C;
            14'd 4700: out = 12'h59C;
            14'd 4701: out = 12'h59C;
            14'd 4702: out = 12'h59C;
            14'd 4703: out = 12'h59C;
            14'd 4704: out = 12'h59C;
            14'd 4705: out = 12'h59D;
            14'd 4706: out = 12'h59D;
            14'd 4707: out = 12'h59D;
            14'd 4708: out = 12'h59D;
            14'd 4709: out = 12'h59D;
            14'd 4710: out = 12'h59D;
            14'd 4711: out = 12'h59D;
            14'd 4712: out = 12'h59D;
            14'd 4713: out = 12'h59E;
            14'd 4714: out = 12'h59E;
            14'd 4715: out = 12'h59E;
            14'd 4716: out = 12'h59E;
            14'd 4717: out = 12'h59E;
            14'd 4718: out = 12'h59E;
            14'd 4719: out = 12'h59E;
            14'd 4720: out = 12'h59E;
            14'd 4721: out = 12'h59E;
            14'd 4722: out = 12'h59F;
            14'd 4723: out = 12'h59F;
            14'd 4724: out = 12'h59F;
            14'd 4725: out = 12'h59F;
            14'd 4726: out = 12'h59F;
            14'd 4727: out = 12'h59F;
            14'd 4728: out = 12'h59F;
            14'd 4729: out = 12'h59F;
            14'd 4730: out = 12'h5A0;
            14'd 4731: out = 12'h5A0;
            14'd 4732: out = 12'h5A0;
            14'd 4733: out = 12'h5A0;
            14'd 4734: out = 12'h5A0;
            14'd 4735: out = 12'h5A0;
            14'd 4736: out = 12'h5A0;
            14'd 4737: out = 12'h5A0;
            14'd 4738: out = 12'h5A1;
            14'd 4739: out = 12'h5A1;
            14'd 4740: out = 12'h5A1;
            14'd 4741: out = 12'h5A1;
            14'd 4742: out = 12'h5A1;
            14'd 4743: out = 12'h5A1;
            14'd 4744: out = 12'h5A1;
            14'd 4745: out = 12'h5A1;
            14'd 4746: out = 12'h5A2;
            14'd 4747: out = 12'h5A2;
            14'd 4748: out = 12'h5A2;
            14'd 4749: out = 12'h5A2;
            14'd 4750: out = 12'h5A2;
            14'd 4751: out = 12'h5A2;
            14'd 4752: out = 12'h5A2;
            14'd 4753: out = 12'h5A2;
            14'd 4754: out = 12'h5A3;
            14'd 4755: out = 12'h5A3;
            14'd 4756: out = 12'h5A3;
            14'd 4757: out = 12'h5A3;
            14'd 4758: out = 12'h5A3;
            14'd 4759: out = 12'h5A3;
            14'd 4760: out = 12'h5A3;
            14'd 4761: out = 12'h5A3;
            14'd 4762: out = 12'h5A4;
            14'd 4763: out = 12'h5A4;
            14'd 4764: out = 12'h5A4;
            14'd 4765: out = 12'h5A4;
            14'd 4766: out = 12'h5A4;
            14'd 4767: out = 12'h5A4;
            14'd 4768: out = 12'h5A4;
            14'd 4769: out = 12'h5A4;
            14'd 4770: out = 12'h5A5;
            14'd 4771: out = 12'h5A5;
            14'd 4772: out = 12'h5A5;
            14'd 4773: out = 12'h5A5;
            14'd 4774: out = 12'h5A5;
            14'd 4775: out = 12'h5A5;
            14'd 4776: out = 12'h5A5;
            14'd 4777: out = 12'h5A5;
            14'd 4778: out = 12'h5A6;
            14'd 4779: out = 12'h5A6;
            14'd 4780: out = 12'h5A6;
            14'd 4781: out = 12'h5A6;
            14'd 4782: out = 12'h5A6;
            14'd 4783: out = 12'h5A6;
            14'd 4784: out = 12'h5A6;
            14'd 4785: out = 12'h5A6;
            14'd 4786: out = 12'h5A7;
            14'd 4787: out = 12'h5A7;
            14'd 4788: out = 12'h5A7;
            14'd 4789: out = 12'h5A7;
            14'd 4790: out = 12'h5A7;
            14'd 4791: out = 12'h5A7;
            14'd 4792: out = 12'h5A7;
            14'd 4793: out = 12'h5A7;
            14'd 4794: out = 12'h5A8;
            14'd 4795: out = 12'h5A8;
            14'd 4796: out = 12'h5A8;
            14'd 4797: out = 12'h5A8;
            14'd 4798: out = 12'h5A8;
            14'd 4799: out = 12'h5A8;
            14'd 4800: out = 12'h5A8;
            14'd 4801: out = 12'h5A8;
            14'd 4802: out = 12'h5A9;
            14'd 4803: out = 12'h5A9;
            14'd 4804: out = 12'h5A9;
            14'd 4805: out = 12'h5A9;
            14'd 4806: out = 12'h5A9;
            14'd 4807: out = 12'h5A9;
            14'd 4808: out = 12'h5A9;
            14'd 4809: out = 12'h5A9;
            14'd 4810: out = 12'h5AA;
            14'd 4811: out = 12'h5AA;
            14'd 4812: out = 12'h5AA;
            14'd 4813: out = 12'h5AA;
            14'd 4814: out = 12'h5AA;
            14'd 4815: out = 12'h5AA;
            14'd 4816: out = 12'h5AA;
            14'd 4817: out = 12'h5AA;
            14'd 4818: out = 12'h5AB;
            14'd 4819: out = 12'h5AB;
            14'd 4820: out = 12'h5AB;
            14'd 4821: out = 12'h5AB;
            14'd 4822: out = 12'h5AB;
            14'd 4823: out = 12'h5AB;
            14'd 4824: out = 12'h5AB;
            14'd 4825: out = 12'h5AB;
            14'd 4826: out = 12'h5AC;
            14'd 4827: out = 12'h5AC;
            14'd 4828: out = 12'h5AC;
            14'd 4829: out = 12'h5AC;
            14'd 4830: out = 12'h5AC;
            14'd 4831: out = 12'h5AC;
            14'd 4832: out = 12'h5AC;
            14'd 4833: out = 12'h5AC;
            14'd 4834: out = 12'h5AD;
            14'd 4835: out = 12'h5AD;
            14'd 4836: out = 12'h5AD;
            14'd 4837: out = 12'h5AD;
            14'd 4838: out = 12'h5AD;
            14'd 4839: out = 12'h5AD;
            14'd 4840: out = 12'h5AD;
            14'd 4841: out = 12'h5AD;
            14'd 4842: out = 12'h5AE;
            14'd 4843: out = 12'h5AE;
            14'd 4844: out = 12'h5AE;
            14'd 4845: out = 12'h5AE;
            14'd 4846: out = 12'h5AE;
            14'd 4847: out = 12'h5AE;
            14'd 4848: out = 12'h5AE;
            14'd 4849: out = 12'h5AE;
            14'd 4850: out = 12'h5AF;
            14'd 4851: out = 12'h5AF;
            14'd 4852: out = 12'h5AF;
            14'd 4853: out = 12'h5AF;
            14'd 4854: out = 12'h5AF;
            14'd 4855: out = 12'h5AF;
            14'd 4856: out = 12'h5AF;
            14'd 4857: out = 12'h5AF;
            14'd 4858: out = 12'h5B0;
            14'd 4859: out = 12'h5B0;
            14'd 4860: out = 12'h5B0;
            14'd 4861: out = 12'h5B0;
            14'd 4862: out = 12'h5B0;
            14'd 4863: out = 12'h5B0;
            14'd 4864: out = 12'h5B0;
            14'd 4865: out = 12'h5B0;
            14'd 4866: out = 12'h5B1;
            14'd 4867: out = 12'h5B1;
            14'd 4868: out = 12'h5B1;
            14'd 4869: out = 12'h5B1;
            14'd 4870: out = 12'h5B1;
            14'd 4871: out = 12'h5B1;
            14'd 4872: out = 12'h5B1;
            14'd 4873: out = 12'h5B1;
            14'd 4874: out = 12'h5B2;
            14'd 4875: out = 12'h5B2;
            14'd 4876: out = 12'h5B2;
            14'd 4877: out = 12'h5B2;
            14'd 4878: out = 12'h5B2;
            14'd 4879: out = 12'h5B2;
            14'd 4880: out = 12'h5B2;
            14'd 4881: out = 12'h5B3;
            14'd 4882: out = 12'h5B3;
            14'd 4883: out = 12'h5B3;
            14'd 4884: out = 12'h5B3;
            14'd 4885: out = 12'h5B3;
            14'd 4886: out = 12'h5B3;
            14'd 4887: out = 12'h5B3;
            14'd 4888: out = 12'h5B3;
            14'd 4889: out = 12'h5B4;
            14'd 4890: out = 12'h5B4;
            14'd 4891: out = 12'h5B4;
            14'd 4892: out = 12'h5B4;
            14'd 4893: out = 12'h5B4;
            14'd 4894: out = 12'h5B4;
            14'd 4895: out = 12'h5B4;
            14'd 4896: out = 12'h5B4;
            14'd 4897: out = 12'h5B5;
            14'd 4898: out = 12'h5B5;
            14'd 4899: out = 12'h5B5;
            14'd 4900: out = 12'h5B5;
            14'd 4901: out = 12'h5B5;
            14'd 4902: out = 12'h5B5;
            14'd 4903: out = 12'h5B5;
            14'd 4904: out = 12'h5B5;
            14'd 4905: out = 12'h5B6;
            14'd 4906: out = 12'h5B6;
            14'd 4907: out = 12'h5B6;
            14'd 4908: out = 12'h5B6;
            14'd 4909: out = 12'h5B6;
            14'd 4910: out = 12'h5B6;
            14'd 4911: out = 12'h5B6;
            14'd 4912: out = 12'h5B6;
            14'd 4913: out = 12'h5B7;
            14'd 4914: out = 12'h5B7;
            14'd 4915: out = 12'h5B7;
            14'd 4916: out = 12'h5B7;
            14'd 4917: out = 12'h5B7;
            14'd 4918: out = 12'h5B7;
            14'd 4919: out = 12'h5B7;
            14'd 4920: out = 12'h5B7;
            14'd 4921: out = 12'h5B8;
            14'd 4922: out = 12'h5B8;
            14'd 4923: out = 12'h5B8;
            14'd 4924: out = 12'h5B8;
            14'd 4925: out = 12'h5B8;
            14'd 4926: out = 12'h5B8;
            14'd 4927: out = 12'h5B8;
            14'd 4928: out = 12'h5B8;
            14'd 4929: out = 12'h5B9;
            14'd 4930: out = 12'h5B9;
            14'd 4931: out = 12'h5B9;
            14'd 4932: out = 12'h5B9;
            14'd 4933: out = 12'h5B9;
            14'd 4934: out = 12'h5B9;
            14'd 4935: out = 12'h5B9;
            14'd 4936: out = 12'h5BA;
            14'd 4937: out = 12'h5BA;
            14'd 4938: out = 12'h5BA;
            14'd 4939: out = 12'h5BA;
            14'd 4940: out = 12'h5BA;
            14'd 4941: out = 12'h5BA;
            14'd 4942: out = 12'h5BA;
            14'd 4943: out = 12'h5BA;
            14'd 4944: out = 12'h5BB;
            14'd 4945: out = 12'h5BB;
            14'd 4946: out = 12'h5BB;
            14'd 4947: out = 12'h5BB;
            14'd 4948: out = 12'h5BB;
            14'd 4949: out = 12'h5BB;
            14'd 4950: out = 12'h5BB;
            14'd 4951: out = 12'h5BB;
            14'd 4952: out = 12'h5BC;
            14'd 4953: out = 12'h5BC;
            14'd 4954: out = 12'h5BC;
            14'd 4955: out = 12'h5BC;
            14'd 4956: out = 12'h5BC;
            14'd 4957: out = 12'h5BC;
            14'd 4958: out = 12'h5BC;
            14'd 4959: out = 12'h5BC;
            14'd 4960: out = 12'h5BD;
            14'd 4961: out = 12'h5BD;
            14'd 4962: out = 12'h5BD;
            14'd 4963: out = 12'h5BD;
            14'd 4964: out = 12'h5BD;
            14'd 4965: out = 12'h5BD;
            14'd 4966: out = 12'h5BD;
            14'd 4967: out = 12'h5BD;
            14'd 4968: out = 12'h5BE;
            14'd 4969: out = 12'h5BE;
            14'd 4970: out = 12'h5BE;
            14'd 4971: out = 12'h5BE;
            14'd 4972: out = 12'h5BE;
            14'd 4973: out = 12'h5BE;
            14'd 4974: out = 12'h5BE;
            14'd 4975: out = 12'h5BF;
            14'd 4976: out = 12'h5BF;
            14'd 4977: out = 12'h5BF;
            14'd 4978: out = 12'h5BF;
            14'd 4979: out = 12'h5BF;
            14'd 4980: out = 12'h5BF;
            14'd 4981: out = 12'h5BF;
            14'd 4982: out = 12'h5BF;
            14'd 4983: out = 12'h5C0;
            14'd 4984: out = 12'h5C0;
            14'd 4985: out = 12'h5C0;
            14'd 4986: out = 12'h5C0;
            14'd 4987: out = 12'h5C0;
            14'd 4988: out = 12'h5C0;
            14'd 4989: out = 12'h5C0;
            14'd 4990: out = 12'h5C0;
            14'd 4991: out = 12'h5C1;
            14'd 4992: out = 12'h5C1;
            14'd 4993: out = 12'h5C1;
            14'd 4994: out = 12'h5C1;
            14'd 4995: out = 12'h5C1;
            14'd 4996: out = 12'h5C1;
            14'd 4997: out = 12'h5C1;
            14'd 4998: out = 12'h5C1;
            14'd 4999: out = 12'h5C2;
            14'd 5000: out = 12'h5C2;
            14'd 5001: out = 12'h5C2;
            14'd 5002: out = 12'h5C2;
            14'd 5003: out = 12'h5C2;
            14'd 5004: out = 12'h5C2;
            14'd 5005: out = 12'h5C2;
            14'd 5006: out = 12'h5C3;
            14'd 5007: out = 12'h5C3;
            14'd 5008: out = 12'h5C3;
            14'd 5009: out = 12'h5C3;
            14'd 5010: out = 12'h5C3;
            14'd 5011: out = 12'h5C3;
            14'd 5012: out = 12'h5C3;
            14'd 5013: out = 12'h5C3;
            14'd 5014: out = 12'h5C4;
            14'd 5015: out = 12'h5C4;
            14'd 5016: out = 12'h5C4;
            14'd 5017: out = 12'h5C4;
            14'd 5018: out = 12'h5C4;
            14'd 5019: out = 12'h5C4;
            14'd 5020: out = 12'h5C4;
            14'd 5021: out = 12'h5C4;
            14'd 5022: out = 12'h5C5;
            14'd 5023: out = 12'h5C5;
            14'd 5024: out = 12'h5C5;
            14'd 5025: out = 12'h5C5;
            14'd 5026: out = 12'h5C5;
            14'd 5027: out = 12'h5C5;
            14'd 5028: out = 12'h5C5;
            14'd 5029: out = 12'h5C6;
            14'd 5030: out = 12'h5C6;
            14'd 5031: out = 12'h5C6;
            14'd 5032: out = 12'h5C6;
            14'd 5033: out = 12'h5C6;
            14'd 5034: out = 12'h5C6;
            14'd 5035: out = 12'h5C6;
            14'd 5036: out = 12'h5C6;
            14'd 5037: out = 12'h5C7;
            14'd 5038: out = 12'h5C7;
            14'd 5039: out = 12'h5C7;
            14'd 5040: out = 12'h5C7;
            14'd 5041: out = 12'h5C7;
            14'd 5042: out = 12'h5C7;
            14'd 5043: out = 12'h5C7;
            14'd 5044: out = 12'h5C7;
            14'd 5045: out = 12'h5C8;
            14'd 5046: out = 12'h5C8;
            14'd 5047: out = 12'h5C8;
            14'd 5048: out = 12'h5C8;
            14'd 5049: out = 12'h5C8;
            14'd 5050: out = 12'h5C8;
            14'd 5051: out = 12'h5C8;
            14'd 5052: out = 12'h5C9;
            14'd 5053: out = 12'h5C9;
            14'd 5054: out = 12'h5C9;
            14'd 5055: out = 12'h5C9;
            14'd 5056: out = 12'h5C9;
            14'd 5057: out = 12'h5C9;
            14'd 5058: out = 12'h5C9;
            14'd 5059: out = 12'h5C9;
            14'd 5060: out = 12'h5CA;
            14'd 5061: out = 12'h5CA;
            14'd 5062: out = 12'h5CA;
            14'd 5063: out = 12'h5CA;
            14'd 5064: out = 12'h5CA;
            14'd 5065: out = 12'h5CA;
            14'd 5066: out = 12'h5CA;
            14'd 5067: out = 12'h5CA;
            14'd 5068: out = 12'h5CB;
            14'd 5069: out = 12'h5CB;
            14'd 5070: out = 12'h5CB;
            14'd 5071: out = 12'h5CB;
            14'd 5072: out = 12'h5CB;
            14'd 5073: out = 12'h5CB;
            14'd 5074: out = 12'h5CB;
            14'd 5075: out = 12'h5CC;
            14'd 5076: out = 12'h5CC;
            14'd 5077: out = 12'h5CC;
            14'd 5078: out = 12'h5CC;
            14'd 5079: out = 12'h5CC;
            14'd 5080: out = 12'h5CC;
            14'd 5081: out = 12'h5CC;
            14'd 5082: out = 12'h5CC;
            14'd 5083: out = 12'h5CD;
            14'd 5084: out = 12'h5CD;
            14'd 5085: out = 12'h5CD;
            14'd 5086: out = 12'h5CD;
            14'd 5087: out = 12'h5CD;
            14'd 5088: out = 12'h5CD;
            14'd 5089: out = 12'h5CD;
            14'd 5090: out = 12'h5CD;
            14'd 5091: out = 12'h5CE;
            14'd 5092: out = 12'h5CE;
            14'd 5093: out = 12'h5CE;
            14'd 5094: out = 12'h5CE;
            14'd 5095: out = 12'h5CE;
            14'd 5096: out = 12'h5CE;
            14'd 5097: out = 12'h5CE;
            14'd 5098: out = 12'h5CF;
            14'd 5099: out = 12'h5CF;
            14'd 5100: out = 12'h5CF;
            14'd 5101: out = 12'h5CF;
            14'd 5102: out = 12'h5CF;
            14'd 5103: out = 12'h5CF;
            14'd 5104: out = 12'h5CF;
            14'd 5105: out = 12'h5CF;
            14'd 5106: out = 12'h5D0;
            14'd 5107: out = 12'h5D0;
            14'd 5108: out = 12'h5D0;
            14'd 5109: out = 12'h5D0;
            14'd 5110: out = 12'h5D0;
            14'd 5111: out = 12'h5D0;
            14'd 5112: out = 12'h5D0;
            14'd 5113: out = 12'h5D1;
            14'd 5114: out = 12'h5D1;
            14'd 5115: out = 12'h5D1;
            14'd 5116: out = 12'h5D1;
            14'd 5117: out = 12'h5D1;
            14'd 5118: out = 12'h5D1;
            14'd 5119: out = 12'h5D1;
            14'd 5120: out = 12'h5D1;
            14'd 5121: out = 12'h5D2;
            14'd 5122: out = 12'h5D2;
            14'd 5123: out = 12'h5D2;
            14'd 5124: out = 12'h5D2;
            14'd 5125: out = 12'h5D2;
            14'd 5126: out = 12'h5D2;
            14'd 5127: out = 12'h5D2;
            14'd 5128: out = 12'h5D3;
            14'd 5129: out = 12'h5D3;
            14'd 5130: out = 12'h5D3;
            14'd 5131: out = 12'h5D3;
            14'd 5132: out = 12'h5D3;
            14'd 5133: out = 12'h5D3;
            14'd 5134: out = 12'h5D3;
            14'd 5135: out = 12'h5D3;
            14'd 5136: out = 12'h5D4;
            14'd 5137: out = 12'h5D4;
            14'd 5138: out = 12'h5D4;
            14'd 5139: out = 12'h5D4;
            14'd 5140: out = 12'h5D4;
            14'd 5141: out = 12'h5D4;
            14'd 5142: out = 12'h5D4;
            14'd 5143: out = 12'h5D5;
            14'd 5144: out = 12'h5D5;
            14'd 5145: out = 12'h5D5;
            14'd 5146: out = 12'h5D5;
            14'd 5147: out = 12'h5D5;
            14'd 5148: out = 12'h5D5;
            14'd 5149: out = 12'h5D5;
            14'd 5150: out = 12'h5D5;
            14'd 5151: out = 12'h5D6;
            14'd 5152: out = 12'h5D6;
            14'd 5153: out = 12'h5D6;
            14'd 5154: out = 12'h5D6;
            14'd 5155: out = 12'h5D6;
            14'd 5156: out = 12'h5D6;
            14'd 5157: out = 12'h5D6;
            14'd 5158: out = 12'h5D6;
            14'd 5159: out = 12'h5D7;
            14'd 5160: out = 12'h5D7;
            14'd 5161: out = 12'h5D7;
            14'd 5162: out = 12'h5D7;
            14'd 5163: out = 12'h5D7;
            14'd 5164: out = 12'h5D7;
            14'd 5165: out = 12'h5D7;
            14'd 5166: out = 12'h5D8;
            14'd 5167: out = 12'h5D8;
            14'd 5168: out = 12'h5D8;
            14'd 5169: out = 12'h5D8;
            14'd 5170: out = 12'h5D8;
            14'd 5171: out = 12'h5D8;
            14'd 5172: out = 12'h5D8;
            14'd 5173: out = 12'h5D8;
            14'd 5174: out = 12'h5D9;
            14'd 5175: out = 12'h5D9;
            14'd 5176: out = 12'h5D9;
            14'd 5177: out = 12'h5D9;
            14'd 5178: out = 12'h5D9;
            14'd 5179: out = 12'h5D9;
            14'd 5180: out = 12'h5D9;
            14'd 5181: out = 12'h5DA;
            14'd 5182: out = 12'h5DA;
            14'd 5183: out = 12'h5DA;
            14'd 5184: out = 12'h5DA;
            14'd 5185: out = 12'h5DA;
            14'd 5186: out = 12'h5DA;
            14'd 5187: out = 12'h5DA;
            14'd 5188: out = 12'h5DB;
            14'd 5189: out = 12'h5DB;
            14'd 5190: out = 12'h5DB;
            14'd 5191: out = 12'h5DB;
            14'd 5192: out = 12'h5DB;
            14'd 5193: out = 12'h5DB;
            14'd 5194: out = 12'h5DB;
            14'd 5195: out = 12'h5DB;
            14'd 5196: out = 12'h5DC;
            14'd 5197: out = 12'h5DC;
            14'd 5198: out = 12'h5DC;
            14'd 5199: out = 12'h5DC;
            14'd 5200: out = 12'h5DC;
            14'd 5201: out = 12'h5DC;
            14'd 5202: out = 12'h5DC;
            14'd 5203: out = 12'h5DD;
            14'd 5204: out = 12'h5DD;
            14'd 5205: out = 12'h5DD;
            14'd 5206: out = 12'h5DD;
            14'd 5207: out = 12'h5DD;
            14'd 5208: out = 12'h5DD;
            14'd 5209: out = 12'h5DD;
            14'd 5210: out = 12'h5DD;
            14'd 5211: out = 12'h5DE;
            14'd 5212: out = 12'h5DE;
            14'd 5213: out = 12'h5DE;
            14'd 5214: out = 12'h5DE;
            14'd 5215: out = 12'h5DE;
            14'd 5216: out = 12'h5DE;
            14'd 5217: out = 12'h5DE;
            14'd 5218: out = 12'h5DF;
            14'd 5219: out = 12'h5DF;
            14'd 5220: out = 12'h5DF;
            14'd 5221: out = 12'h5DF;
            14'd 5222: out = 12'h5DF;
            14'd 5223: out = 12'h5DF;
            14'd 5224: out = 12'h5DF;
            14'd 5225: out = 12'h5DF;
            14'd 5226: out = 12'h5E0;
            14'd 5227: out = 12'h5E0;
            14'd 5228: out = 12'h5E0;
            14'd 5229: out = 12'h5E0;
            14'd 5230: out = 12'h5E0;
            14'd 5231: out = 12'h5E0;
            14'd 5232: out = 12'h5E0;
            14'd 5233: out = 12'h5E1;
            14'd 5234: out = 12'h5E1;
            14'd 5235: out = 12'h5E1;
            14'd 5236: out = 12'h5E1;
            14'd 5237: out = 12'h5E1;
            14'd 5238: out = 12'h5E1;
            14'd 5239: out = 12'h5E1;
            14'd 5240: out = 12'h5E1;
            14'd 5241: out = 12'h5E2;
            14'd 5242: out = 12'h5E2;
            14'd 5243: out = 12'h5E2;
            14'd 5244: out = 12'h5E2;
            14'd 5245: out = 12'h5E2;
            14'd 5246: out = 12'h5E2;
            14'd 5247: out = 12'h5E2;
            14'd 5248: out = 12'h5E3;
            14'd 5249: out = 12'h5E3;
            14'd 5250: out = 12'h5E3;
            14'd 5251: out = 12'h5E3;
            14'd 5252: out = 12'h5E3;
            14'd 5253: out = 12'h5E3;
            14'd 5254: out = 12'h5E3;
            14'd 5255: out = 12'h5E4;
            14'd 5256: out = 12'h5E4;
            14'd 5257: out = 12'h5E4;
            14'd 5258: out = 12'h5E4;
            14'd 5259: out = 12'h5E4;
            14'd 5260: out = 12'h5E4;
            14'd 5261: out = 12'h5E4;
            14'd 5262: out = 12'h5E4;
            14'd 5263: out = 12'h5E5;
            14'd 5264: out = 12'h5E5;
            14'd 5265: out = 12'h5E5;
            14'd 5266: out = 12'h5E5;
            14'd 5267: out = 12'h5E5;
            14'd 5268: out = 12'h5E5;
            14'd 5269: out = 12'h5E5;
            14'd 5270: out = 12'h5E6;
            14'd 5271: out = 12'h5E6;
            14'd 5272: out = 12'h5E6;
            14'd 5273: out = 12'h5E6;
            14'd 5274: out = 12'h5E6;
            14'd 5275: out = 12'h5E6;
            14'd 5276: out = 12'h5E6;
            14'd 5277: out = 12'h5E7;
            14'd 5278: out = 12'h5E7;
            14'd 5279: out = 12'h5E7;
            14'd 5280: out = 12'h5E7;
            14'd 5281: out = 12'h5E7;
            14'd 5282: out = 12'h5E7;
            14'd 5283: out = 12'h5E7;
            14'd 5284: out = 12'h5E7;
            14'd 5285: out = 12'h5E8;
            14'd 5286: out = 12'h5E8;
            14'd 5287: out = 12'h5E8;
            14'd 5288: out = 12'h5E8;
            14'd 5289: out = 12'h5E8;
            14'd 5290: out = 12'h5E8;
            14'd 5291: out = 12'h5E8;
            14'd 5292: out = 12'h5E9;
            14'd 5293: out = 12'h5E9;
            14'd 5294: out = 12'h5E9;
            14'd 5295: out = 12'h5E9;
            14'd 5296: out = 12'h5E9;
            14'd 5297: out = 12'h5E9;
            14'd 5298: out = 12'h5E9;
            14'd 5299: out = 12'h5EA;
            14'd 5300: out = 12'h5EA;
            14'd 5301: out = 12'h5EA;
            14'd 5302: out = 12'h5EA;
            14'd 5303: out = 12'h5EA;
            14'd 5304: out = 12'h5EA;
            14'd 5305: out = 12'h5EA;
            14'd 5306: out = 12'h5EA;
            14'd 5307: out = 12'h5EB;
            14'd 5308: out = 12'h5EB;
            14'd 5309: out = 12'h5EB;
            14'd 5310: out = 12'h5EB;
            14'd 5311: out = 12'h5EB;
            14'd 5312: out = 12'h5EB;
            14'd 5313: out = 12'h5EB;
            14'd 5314: out = 12'h5EC;
            14'd 5315: out = 12'h5EC;
            14'd 5316: out = 12'h5EC;
            14'd 5317: out = 12'h5EC;
            14'd 5318: out = 12'h5EC;
            14'd 5319: out = 12'h5EC;
            14'd 5320: out = 12'h5EC;
            14'd 5321: out = 12'h5ED;
            14'd 5322: out = 12'h5ED;
            14'd 5323: out = 12'h5ED;
            14'd 5324: out = 12'h5ED;
            14'd 5325: out = 12'h5ED;
            14'd 5326: out = 12'h5ED;
            14'd 5327: out = 12'h5ED;
            14'd 5328: out = 12'h5ED;
            14'd 5329: out = 12'h5EE;
            14'd 5330: out = 12'h5EE;
            14'd 5331: out = 12'h5EE;
            14'd 5332: out = 12'h5EE;
            14'd 5333: out = 12'h5EE;
            14'd 5334: out = 12'h5EE;
            14'd 5335: out = 12'h5EE;
            14'd 5336: out = 12'h5EF;
            14'd 5337: out = 12'h5EF;
            14'd 5338: out = 12'h5EF;
            14'd 5339: out = 12'h5EF;
            14'd 5340: out = 12'h5EF;
            14'd 5341: out = 12'h5EF;
            14'd 5342: out = 12'h5EF;
            14'd 5343: out = 12'h5F0;
            14'd 5344: out = 12'h5F0;
            14'd 5345: out = 12'h5F0;
            14'd 5346: out = 12'h5F0;
            14'd 5347: out = 12'h5F0;
            14'd 5348: out = 12'h5F0;
            14'd 5349: out = 12'h5F0;
            14'd 5350: out = 12'h5F1;
            14'd 5351: out = 12'h5F1;
            14'd 5352: out = 12'h5F1;
            14'd 5353: out = 12'h5F1;
            14'd 5354: out = 12'h5F1;
            14'd 5355: out = 12'h5F1;
            14'd 5356: out = 12'h5F1;
            14'd 5357: out = 12'h5F1;
            14'd 5358: out = 12'h5F2;
            14'd 5359: out = 12'h5F2;
            14'd 5360: out = 12'h5F2;
            14'd 5361: out = 12'h5F2;
            14'd 5362: out = 12'h5F2;
            14'd 5363: out = 12'h5F2;
            14'd 5364: out = 12'h5F2;
            14'd 5365: out = 12'h5F3;
            14'd 5366: out = 12'h5F3;
            14'd 5367: out = 12'h5F3;
            14'd 5368: out = 12'h5F3;
            14'd 5369: out = 12'h5F3;
            14'd 5370: out = 12'h5F3;
            14'd 5371: out = 12'h5F3;
            14'd 5372: out = 12'h5F4;
            14'd 5373: out = 12'h5F4;
            14'd 5374: out = 12'h5F4;
            14'd 5375: out = 12'h5F4;
            14'd 5376: out = 12'h5F4;
            14'd 5377: out = 12'h5F4;
            14'd 5378: out = 12'h5F4;
            14'd 5379: out = 12'h5F5;
            14'd 5380: out = 12'h5F5;
            14'd 5381: out = 12'h5F5;
            14'd 5382: out = 12'h5F5;
            14'd 5383: out = 12'h5F5;
            14'd 5384: out = 12'h5F5;
            14'd 5385: out = 12'h5F5;
            14'd 5386: out = 12'h5F5;
            14'd 5387: out = 12'h5F6;
            14'd 5388: out = 12'h5F6;
            14'd 5389: out = 12'h5F6;
            14'd 5390: out = 12'h5F6;
            14'd 5391: out = 12'h5F6;
            14'd 5392: out = 12'h5F6;
            14'd 5393: out = 12'h5F6;
            14'd 5394: out = 12'h5F7;
            14'd 5395: out = 12'h5F7;
            14'd 5396: out = 12'h5F7;
            14'd 5397: out = 12'h5F7;
            14'd 5398: out = 12'h5F7;
            14'd 5399: out = 12'h5F7;
            14'd 5400: out = 12'h5F7;
            14'd 5401: out = 12'h5F8;
            14'd 5402: out = 12'h5F8;
            14'd 5403: out = 12'h5F8;
            14'd 5404: out = 12'h5F8;
            14'd 5405: out = 12'h5F8;
            14'd 5406: out = 12'h5F8;
            14'd 5407: out = 12'h5F8;
            14'd 5408: out = 12'h5F9;
            14'd 5409: out = 12'h5F9;
            14'd 5410: out = 12'h5F9;
            14'd 5411: out = 12'h5F9;
            14'd 5412: out = 12'h5F9;
            14'd 5413: out = 12'h5F9;
            14'd 5414: out = 12'h5F9;
            14'd 5415: out = 12'h5FA;
            14'd 5416: out = 12'h5FA;
            14'd 5417: out = 12'h5FA;
            14'd 5418: out = 12'h5FA;
            14'd 5419: out = 12'h5FA;
            14'd 5420: out = 12'h5FA;
            14'd 5421: out = 12'h5FA;
            14'd 5422: out = 12'h5FA;
            14'd 5423: out = 12'h5FB;
            14'd 5424: out = 12'h5FB;
            14'd 5425: out = 12'h5FB;
            14'd 5426: out = 12'h5FB;
            14'd 5427: out = 12'h5FB;
            14'd 5428: out = 12'h5FB;
            14'd 5429: out = 12'h5FB;
            14'd 5430: out = 12'h5FC;
            14'd 5431: out = 12'h5FC;
            14'd 5432: out = 12'h5FC;
            14'd 5433: out = 12'h5FC;
            14'd 5434: out = 12'h5FC;
            14'd 5435: out = 12'h5FC;
            14'd 5436: out = 12'h5FC;
            14'd 5437: out = 12'h5FD;
            14'd 5438: out = 12'h5FD;
            14'd 5439: out = 12'h5FD;
            14'd 5440: out = 12'h5FD;
            14'd 5441: out = 12'h5FD;
            14'd 5442: out = 12'h5FD;
            14'd 5443: out = 12'h5FD;
            14'd 5444: out = 12'h5FE;
            14'd 5445: out = 12'h5FE;
            14'd 5446: out = 12'h5FE;
            14'd 5447: out = 12'h5FE;
            14'd 5448: out = 12'h5FE;
            14'd 5449: out = 12'h5FE;
            14'd 5450: out = 12'h5FE;
            14'd 5451: out = 12'h5FF;
            14'd 5452: out = 12'h5FF;
            14'd 5453: out = 12'h5FF;
            14'd 5454: out = 12'h5FF;
            14'd 5455: out = 12'h5FF;
            14'd 5456: out = 12'h5FF;
            14'd 5457: out = 12'h5FF;
            14'd 5458: out = 12'h600;
            14'd 5459: out = 12'h600;
            14'd 5460: out = 12'h600;
            14'd 5461: out = 12'h600;
            14'd 5462: out = 12'h600;
            14'd 5463: out = 12'h600;
            14'd 5464: out = 12'h600;
            14'd 5465: out = 12'h601;
            14'd 5466: out = 12'h601;
            14'd 5467: out = 12'h601;
            14'd 5468: out = 12'h601;
            14'd 5469: out = 12'h601;
            14'd 5470: out = 12'h601;
            14'd 5471: out = 12'h601;
            14'd 5472: out = 12'h602;
            14'd 5473: out = 12'h602;
            14'd 5474: out = 12'h602;
            14'd 5475: out = 12'h602;
            14'd 5476: out = 12'h602;
            14'd 5477: out = 12'h602;
            14'd 5478: out = 12'h602;
            14'd 5479: out = 12'h602;
            14'd 5480: out = 12'h603;
            14'd 5481: out = 12'h603;
            14'd 5482: out = 12'h603;
            14'd 5483: out = 12'h603;
            14'd 5484: out = 12'h603;
            14'd 5485: out = 12'h603;
            14'd 5486: out = 12'h603;
            14'd 5487: out = 12'h604;
            14'd 5488: out = 12'h604;
            14'd 5489: out = 12'h604;
            14'd 5490: out = 12'h604;
            14'd 5491: out = 12'h604;
            14'd 5492: out = 12'h604;
            14'd 5493: out = 12'h604;
            14'd 5494: out = 12'h605;
            14'd 5495: out = 12'h605;
            14'd 5496: out = 12'h605;
            14'd 5497: out = 12'h605;
            14'd 5498: out = 12'h605;
            14'd 5499: out = 12'h605;
            14'd 5500: out = 12'h605;
            14'd 5501: out = 12'h606;
            14'd 5502: out = 12'h606;
            14'd 5503: out = 12'h606;
            14'd 5504: out = 12'h606;
            14'd 5505: out = 12'h606;
            14'd 5506: out = 12'h606;
            14'd 5507: out = 12'h606;
            14'd 5508: out = 12'h607;
            14'd 5509: out = 12'h607;
            14'd 5510: out = 12'h607;
            14'd 5511: out = 12'h607;
            14'd 5512: out = 12'h607;
            14'd 5513: out = 12'h607;
            14'd 5514: out = 12'h607;
            14'd 5515: out = 12'h608;
            14'd 5516: out = 12'h608;
            14'd 5517: out = 12'h608;
            14'd 5518: out = 12'h608;
            14'd 5519: out = 12'h608;
            14'd 5520: out = 12'h608;
            14'd 5521: out = 12'h608;
            14'd 5522: out = 12'h609;
            14'd 5523: out = 12'h609;
            14'd 5524: out = 12'h609;
            14'd 5525: out = 12'h609;
            14'd 5526: out = 12'h609;
            14'd 5527: out = 12'h609;
            14'd 5528: out = 12'h609;
            14'd 5529: out = 12'h60A;
            14'd 5530: out = 12'h60A;
            14'd 5531: out = 12'h60A;
            14'd 5532: out = 12'h60A;
            14'd 5533: out = 12'h60A;
            14'd 5534: out = 12'h60A;
            14'd 5535: out = 12'h60A;
            14'd 5536: out = 12'h60B;
            14'd 5537: out = 12'h60B;
            14'd 5538: out = 12'h60B;
            14'd 5539: out = 12'h60B;
            14'd 5540: out = 12'h60B;
            14'd 5541: out = 12'h60B;
            14'd 5542: out = 12'h60B;
            14'd 5543: out = 12'h60C;
            14'd 5544: out = 12'h60C;
            14'd 5545: out = 12'h60C;
            14'd 5546: out = 12'h60C;
            14'd 5547: out = 12'h60C;
            14'd 5548: out = 12'h60C;
            14'd 5549: out = 12'h60C;
            14'd 5550: out = 12'h60D;
            14'd 5551: out = 12'h60D;
            14'd 5552: out = 12'h60D;
            14'd 5553: out = 12'h60D;
            14'd 5554: out = 12'h60D;
            14'd 5555: out = 12'h60D;
            14'd 5556: out = 12'h60D;
            14'd 5557: out = 12'h60E;
            14'd 5558: out = 12'h60E;
            14'd 5559: out = 12'h60E;
            14'd 5560: out = 12'h60E;
            14'd 5561: out = 12'h60E;
            14'd 5562: out = 12'h60E;
            14'd 5563: out = 12'h60E;
            14'd 5564: out = 12'h60F;
            14'd 5565: out = 12'h60F;
            14'd 5566: out = 12'h60F;
            14'd 5567: out = 12'h60F;
            14'd 5568: out = 12'h60F;
            14'd 5569: out = 12'h60F;
            14'd 5570: out = 12'h60F;
            14'd 5571: out = 12'h610;
            14'd 5572: out = 12'h610;
            14'd 5573: out = 12'h610;
            14'd 5574: out = 12'h610;
            14'd 5575: out = 12'h610;
            14'd 5576: out = 12'h610;
            14'd 5577: out = 12'h610;
            14'd 5578: out = 12'h611;
            14'd 5579: out = 12'h611;
            14'd 5580: out = 12'h611;
            14'd 5581: out = 12'h611;
            14'd 5582: out = 12'h611;
            14'd 5583: out = 12'h611;
            14'd 5584: out = 12'h611;
            14'd 5585: out = 12'h612;
            14'd 5586: out = 12'h612;
            14'd 5587: out = 12'h612;
            14'd 5588: out = 12'h612;
            14'd 5589: out = 12'h612;
            14'd 5590: out = 12'h612;
            14'd 5591: out = 12'h612;
            14'd 5592: out = 12'h613;
            14'd 5593: out = 12'h613;
            14'd 5594: out = 12'h613;
            14'd 5595: out = 12'h613;
            14'd 5596: out = 12'h613;
            14'd 5597: out = 12'h613;
            14'd 5598: out = 12'h613;
            14'd 5599: out = 12'h614;
            14'd 5600: out = 12'h614;
            14'd 5601: out = 12'h614;
            14'd 5602: out = 12'h614;
            14'd 5603: out = 12'h614;
            14'd 5604: out = 12'h614;
            14'd 5605: out = 12'h614;
            14'd 5606: out = 12'h615;
            14'd 5607: out = 12'h615;
            14'd 5608: out = 12'h615;
            14'd 5609: out = 12'h615;
            14'd 5610: out = 12'h615;
            14'd 5611: out = 12'h615;
            14'd 5612: out = 12'h615;
            14'd 5613: out = 12'h616;
            14'd 5614: out = 12'h616;
            14'd 5615: out = 12'h616;
            14'd 5616: out = 12'h616;
            14'd 5617: out = 12'h616;
            14'd 5618: out = 12'h616;
            14'd 5619: out = 12'h616;
            14'd 5620: out = 12'h617;
            14'd 5621: out = 12'h617;
            14'd 5622: out = 12'h617;
            14'd 5623: out = 12'h617;
            14'd 5624: out = 12'h617;
            14'd 5625: out = 12'h617;
            14'd 5626: out = 12'h618;
            14'd 5627: out = 12'h618;
            14'd 5628: out = 12'h618;
            14'd 5629: out = 12'h618;
            14'd 5630: out = 12'h618;
            14'd 5631: out = 12'h618;
            14'd 5632: out = 12'h618;
            14'd 5633: out = 12'h619;
            14'd 5634: out = 12'h619;
            14'd 5635: out = 12'h619;
            14'd 5636: out = 12'h619;
            14'd 5637: out = 12'h619;
            14'd 5638: out = 12'h619;
            14'd 5639: out = 12'h619;
            14'd 5640: out = 12'h61A;
            14'd 5641: out = 12'h61A;
            14'd 5642: out = 12'h61A;
            14'd 5643: out = 12'h61A;
            14'd 5644: out = 12'h61A;
            14'd 5645: out = 12'h61A;
            14'd 5646: out = 12'h61A;
            14'd 5647: out = 12'h61B;
            14'd 5648: out = 12'h61B;
            14'd 5649: out = 12'h61B;
            14'd 5650: out = 12'h61B;
            14'd 5651: out = 12'h61B;
            14'd 5652: out = 12'h61B;
            14'd 5653: out = 12'h61B;
            14'd 5654: out = 12'h61C;
            14'd 5655: out = 12'h61C;
            14'd 5656: out = 12'h61C;
            14'd 5657: out = 12'h61C;
            14'd 5658: out = 12'h61C;
            14'd 5659: out = 12'h61C;
            14'd 5660: out = 12'h61C;
            14'd 5661: out = 12'h61D;
            14'd 5662: out = 12'h61D;
            14'd 5663: out = 12'h61D;
            14'd 5664: out = 12'h61D;
            14'd 5665: out = 12'h61D;
            14'd 5666: out = 12'h61D;
            14'd 5667: out = 12'h61D;
            14'd 5668: out = 12'h61E;
            14'd 5669: out = 12'h61E;
            14'd 5670: out = 12'h61E;
            14'd 5671: out = 12'h61E;
            14'd 5672: out = 12'h61E;
            14'd 5673: out = 12'h61E;
            14'd 5674: out = 12'h61F;
            14'd 5675: out = 12'h61F;
            14'd 5676: out = 12'h61F;
            14'd 5677: out = 12'h61F;
            14'd 5678: out = 12'h61F;
            14'd 5679: out = 12'h61F;
            14'd 5680: out = 12'h61F;
            14'd 5681: out = 12'h620;
            14'd 5682: out = 12'h620;
            14'd 5683: out = 12'h620;
            14'd 5684: out = 12'h620;
            14'd 5685: out = 12'h620;
            14'd 5686: out = 12'h620;
            14'd 5687: out = 12'h620;
            14'd 5688: out = 12'h621;
            14'd 5689: out = 12'h621;
            14'd 5690: out = 12'h621;
            14'd 5691: out = 12'h621;
            14'd 5692: out = 12'h621;
            14'd 5693: out = 12'h621;
            14'd 5694: out = 12'h621;
            14'd 5695: out = 12'h622;
            14'd 5696: out = 12'h622;
            14'd 5697: out = 12'h622;
            14'd 5698: out = 12'h622;
            14'd 5699: out = 12'h622;
            14'd 5700: out = 12'h622;
            14'd 5701: out = 12'h622;
            14'd 5702: out = 12'h623;
            14'd 5703: out = 12'h623;
            14'd 5704: out = 12'h623;
            14'd 5705: out = 12'h623;
            14'd 5706: out = 12'h623;
            14'd 5707: out = 12'h623;
            14'd 5708: out = 12'h623;
            14'd 5709: out = 12'h624;
            14'd 5710: out = 12'h624;
            14'd 5711: out = 12'h624;
            14'd 5712: out = 12'h624;
            14'd 5713: out = 12'h624;
            14'd 5714: out = 12'h624;
            14'd 5715: out = 12'h625;
            14'd 5716: out = 12'h625;
            14'd 5717: out = 12'h625;
            14'd 5718: out = 12'h625;
            14'd 5719: out = 12'h625;
            14'd 5720: out = 12'h625;
            14'd 5721: out = 12'h625;
            14'd 5722: out = 12'h626;
            14'd 5723: out = 12'h626;
            14'd 5724: out = 12'h626;
            14'd 5725: out = 12'h626;
            14'd 5726: out = 12'h626;
            14'd 5727: out = 12'h626;
            14'd 5728: out = 12'h626;
            14'd 5729: out = 12'h627;
            14'd 5730: out = 12'h627;
            14'd 5731: out = 12'h627;
            14'd 5732: out = 12'h627;
            14'd 5733: out = 12'h627;
            14'd 5734: out = 12'h627;
            14'd 5735: out = 12'h627;
            14'd 5736: out = 12'h628;
            14'd 5737: out = 12'h628;
            14'd 5738: out = 12'h628;
            14'd 5739: out = 12'h628;
            14'd 5740: out = 12'h628;
            14'd 5741: out = 12'h628;
            14'd 5742: out = 12'h629;
            14'd 5743: out = 12'h629;
            14'd 5744: out = 12'h629;
            14'd 5745: out = 12'h629;
            14'd 5746: out = 12'h629;
            14'd 5747: out = 12'h629;
            14'd 5748: out = 12'h629;
            14'd 5749: out = 12'h62A;
            14'd 5750: out = 12'h62A;
            14'd 5751: out = 12'h62A;
            14'd 5752: out = 12'h62A;
            14'd 5753: out = 12'h62A;
            14'd 5754: out = 12'h62A;
            14'd 5755: out = 12'h62A;
            14'd 5756: out = 12'h62B;
            14'd 5757: out = 12'h62B;
            14'd 5758: out = 12'h62B;
            14'd 5759: out = 12'h62B;
            14'd 5760: out = 12'h62B;
            14'd 5761: out = 12'h62B;
            14'd 5762: out = 12'h62B;
            14'd 5763: out = 12'h62C;
            14'd 5764: out = 12'h62C;
            14'd 5765: out = 12'h62C;
            14'd 5766: out = 12'h62C;
            14'd 5767: out = 12'h62C;
            14'd 5768: out = 12'h62C;
            14'd 5769: out = 12'h62D;
            14'd 5770: out = 12'h62D;
            14'd 5771: out = 12'h62D;
            14'd 5772: out = 12'h62D;
            14'd 5773: out = 12'h62D;
            14'd 5774: out = 12'h62D;
            14'd 5775: out = 12'h62D;
            14'd 5776: out = 12'h62E;
            14'd 5777: out = 12'h62E;
            14'd 5778: out = 12'h62E;
            14'd 5779: out = 12'h62E;
            14'd 5780: out = 12'h62E;
            14'd 5781: out = 12'h62E;
            14'd 5782: out = 12'h62E;
            14'd 5783: out = 12'h62F;
            14'd 5784: out = 12'h62F;
            14'd 5785: out = 12'h62F;
            14'd 5786: out = 12'h62F;
            14'd 5787: out = 12'h62F;
            14'd 5788: out = 12'h62F;
            14'd 5789: out = 12'h630;
            14'd 5790: out = 12'h630;
            14'd 5791: out = 12'h630;
            14'd 5792: out = 12'h630;
            14'd 5793: out = 12'h630;
            14'd 5794: out = 12'h630;
            14'd 5795: out = 12'h630;
            14'd 5796: out = 12'h631;
            14'd 5797: out = 12'h631;
            14'd 5798: out = 12'h631;
            14'd 5799: out = 12'h631;
            14'd 5800: out = 12'h631;
            14'd 5801: out = 12'h631;
            14'd 5802: out = 12'h631;
            14'd 5803: out = 12'h632;
            14'd 5804: out = 12'h632;
            14'd 5805: out = 12'h632;
            14'd 5806: out = 12'h632;
            14'd 5807: out = 12'h632;
            14'd 5808: out = 12'h632;
            14'd 5809: out = 12'h632;
            14'd 5810: out = 12'h633;
            14'd 5811: out = 12'h633;
            14'd 5812: out = 12'h633;
            14'd 5813: out = 12'h633;
            14'd 5814: out = 12'h633;
            14'd 5815: out = 12'h633;
            14'd 5816: out = 12'h634;
            14'd 5817: out = 12'h634;
            14'd 5818: out = 12'h634;
            14'd 5819: out = 12'h634;
            14'd 5820: out = 12'h634;
            14'd 5821: out = 12'h634;
            14'd 5822: out = 12'h634;
            14'd 5823: out = 12'h635;
            14'd 5824: out = 12'h635;
            14'd 5825: out = 12'h635;
            14'd 5826: out = 12'h635;
            14'd 5827: out = 12'h635;
            14'd 5828: out = 12'h635;
            14'd 5829: out = 12'h636;
            14'd 5830: out = 12'h636;
            14'd 5831: out = 12'h636;
            14'd 5832: out = 12'h636;
            14'd 5833: out = 12'h636;
            14'd 5834: out = 12'h636;
            14'd 5835: out = 12'h636;
            14'd 5836: out = 12'h637;
            14'd 5837: out = 12'h637;
            14'd 5838: out = 12'h637;
            14'd 5839: out = 12'h637;
            14'd 5840: out = 12'h637;
            14'd 5841: out = 12'h637;
            14'd 5842: out = 12'h637;
            14'd 5843: out = 12'h638;
            14'd 5844: out = 12'h638;
            14'd 5845: out = 12'h638;
            14'd 5846: out = 12'h638;
            14'd 5847: out = 12'h638;
            14'd 5848: out = 12'h638;
            14'd 5849: out = 12'h639;
            14'd 5850: out = 12'h639;
            14'd 5851: out = 12'h639;
            14'd 5852: out = 12'h639;
            14'd 5853: out = 12'h639;
            14'd 5854: out = 12'h639;
            14'd 5855: out = 12'h639;
            14'd 5856: out = 12'h63A;
            14'd 5857: out = 12'h63A;
            14'd 5858: out = 12'h63A;
            14'd 5859: out = 12'h63A;
            14'd 5860: out = 12'h63A;
            14'd 5861: out = 12'h63A;
            14'd 5862: out = 12'h63A;
            14'd 5863: out = 12'h63B;
            14'd 5864: out = 12'h63B;
            14'd 5865: out = 12'h63B;
            14'd 5866: out = 12'h63B;
            14'd 5867: out = 12'h63B;
            14'd 5868: out = 12'h63B;
            14'd 5869: out = 12'h63C;
            14'd 5870: out = 12'h63C;
            14'd 5871: out = 12'h63C;
            14'd 5872: out = 12'h63C;
            14'd 5873: out = 12'h63C;
            14'd 5874: out = 12'h63C;
            14'd 5875: out = 12'h63C;
            14'd 5876: out = 12'h63D;
            14'd 5877: out = 12'h63D;
            14'd 5878: out = 12'h63D;
            14'd 5879: out = 12'h63D;
            14'd 5880: out = 12'h63D;
            14'd 5881: out = 12'h63D;
            14'd 5882: out = 12'h63E;
            14'd 5883: out = 12'h63E;
            14'd 5884: out = 12'h63E;
            14'd 5885: out = 12'h63E;
            14'd 5886: out = 12'h63E;
            14'd 5887: out = 12'h63E;
            14'd 5888: out = 12'h63E;
            14'd 5889: out = 12'h63F;
            14'd 5890: out = 12'h63F;
            14'd 5891: out = 12'h63F;
            14'd 5892: out = 12'h63F;
            14'd 5893: out = 12'h63F;
            14'd 5894: out = 12'h63F;
            14'd 5895: out = 12'h640;
            14'd 5896: out = 12'h640;
            14'd 5897: out = 12'h640;
            14'd 5898: out = 12'h640;
            14'd 5899: out = 12'h640;
            14'd 5900: out = 12'h640;
            14'd 5901: out = 12'h640;
            14'd 5902: out = 12'h641;
            14'd 5903: out = 12'h641;
            14'd 5904: out = 12'h641;
            14'd 5905: out = 12'h641;
            14'd 5906: out = 12'h641;
            14'd 5907: out = 12'h641;
            14'd 5908: out = 12'h641;
            14'd 5909: out = 12'h642;
            14'd 5910: out = 12'h642;
            14'd 5911: out = 12'h642;
            14'd 5912: out = 12'h642;
            14'd 5913: out = 12'h642;
            14'd 5914: out = 12'h642;
            14'd 5915: out = 12'h643;
            14'd 5916: out = 12'h643;
            14'd 5917: out = 12'h643;
            14'd 5918: out = 12'h643;
            14'd 5919: out = 12'h643;
            14'd 5920: out = 12'h643;
            14'd 5921: out = 12'h643;
            14'd 5922: out = 12'h644;
            14'd 5923: out = 12'h644;
            14'd 5924: out = 12'h644;
            14'd 5925: out = 12'h644;
            14'd 5926: out = 12'h644;
            14'd 5927: out = 12'h644;
            14'd 5928: out = 12'h645;
            14'd 5929: out = 12'h645;
            14'd 5930: out = 12'h645;
            14'd 5931: out = 12'h645;
            14'd 5932: out = 12'h645;
            14'd 5933: out = 12'h645;
            14'd 5934: out = 12'h645;
            14'd 5935: out = 12'h646;
            14'd 5936: out = 12'h646;
            14'd 5937: out = 12'h646;
            14'd 5938: out = 12'h646;
            14'd 5939: out = 12'h646;
            14'd 5940: out = 12'h646;
            14'd 5941: out = 12'h647;
            14'd 5942: out = 12'h647;
            14'd 5943: out = 12'h647;
            14'd 5944: out = 12'h647;
            14'd 5945: out = 12'h647;
            14'd 5946: out = 12'h647;
            14'd 5947: out = 12'h647;
            14'd 5948: out = 12'h648;
            14'd 5949: out = 12'h648;
            14'd 5950: out = 12'h648;
            14'd 5951: out = 12'h648;
            14'd 5952: out = 12'h648;
            14'd 5953: out = 12'h648;
            14'd 5954: out = 12'h649;
            14'd 5955: out = 12'h649;
            14'd 5956: out = 12'h649;
            14'd 5957: out = 12'h649;
            14'd 5958: out = 12'h649;
            14'd 5959: out = 12'h649;
            14'd 5960: out = 12'h649;
            14'd 5961: out = 12'h64A;
            14'd 5962: out = 12'h64A;
            14'd 5963: out = 12'h64A;
            14'd 5964: out = 12'h64A;
            14'd 5965: out = 12'h64A;
            14'd 5966: out = 12'h64A;
            14'd 5967: out = 12'h64B;
            14'd 5968: out = 12'h64B;
            14'd 5969: out = 12'h64B;
            14'd 5970: out = 12'h64B;
            14'd 5971: out = 12'h64B;
            14'd 5972: out = 12'h64B;
            14'd 5973: out = 12'h64B;
            14'd 5974: out = 12'h64C;
            14'd 5975: out = 12'h64C;
            14'd 5976: out = 12'h64C;
            14'd 5977: out = 12'h64C;
            14'd 5978: out = 12'h64C;
            14'd 5979: out = 12'h64C;
            14'd 5980: out = 12'h64D;
            14'd 5981: out = 12'h64D;
            14'd 5982: out = 12'h64D;
            14'd 5983: out = 12'h64D;
            14'd 5984: out = 12'h64D;
            14'd 5985: out = 12'h64D;
            14'd 5986: out = 12'h64E;
            14'd 5987: out = 12'h64E;
            14'd 5988: out = 12'h64E;
            14'd 5989: out = 12'h64E;
            14'd 5990: out = 12'h64E;
            14'd 5991: out = 12'h64E;
            14'd 5992: out = 12'h64E;
            14'd 5993: out = 12'h64F;
            14'd 5994: out = 12'h64F;
            14'd 5995: out = 12'h64F;
            14'd 5996: out = 12'h64F;
            14'd 5997: out = 12'h64F;
            14'd 5998: out = 12'h64F;
            14'd 5999: out = 12'h650;
            14'd 6000: out = 12'h650;
            14'd 6001: out = 12'h650;
            14'd 6002: out = 12'h650;
            14'd 6003: out = 12'h650;
            14'd 6004: out = 12'h650;
            14'd 6005: out = 12'h650;
            14'd 6006: out = 12'h651;
            14'd 6007: out = 12'h651;
            14'd 6008: out = 12'h651;
            14'd 6009: out = 12'h651;
            14'd 6010: out = 12'h651;
            14'd 6011: out = 12'h651;
            14'd 6012: out = 12'h652;
            14'd 6013: out = 12'h652;
            14'd 6014: out = 12'h652;
            14'd 6015: out = 12'h652;
            14'd 6016: out = 12'h652;
            14'd 6017: out = 12'h652;
            14'd 6018: out = 12'h652;
            14'd 6019: out = 12'h653;
            14'd 6020: out = 12'h653;
            14'd 6021: out = 12'h653;
            14'd 6022: out = 12'h653;
            14'd 6023: out = 12'h653;
            14'd 6024: out = 12'h653;
            14'd 6025: out = 12'h654;
            14'd 6026: out = 12'h654;
            14'd 6027: out = 12'h654;
            14'd 6028: out = 12'h654;
            14'd 6029: out = 12'h654;
            14'd 6030: out = 12'h654;
            14'd 6031: out = 12'h655;
            14'd 6032: out = 12'h655;
            14'd 6033: out = 12'h655;
            14'd 6034: out = 12'h655;
            14'd 6035: out = 12'h655;
            14'd 6036: out = 12'h655;
            14'd 6037: out = 12'h655;
            14'd 6038: out = 12'h656;
            14'd 6039: out = 12'h656;
            14'd 6040: out = 12'h656;
            14'd 6041: out = 12'h656;
            14'd 6042: out = 12'h656;
            14'd 6043: out = 12'h656;
            14'd 6044: out = 12'h657;
            14'd 6045: out = 12'h657;
            14'd 6046: out = 12'h657;
            14'd 6047: out = 12'h657;
            14'd 6048: out = 12'h657;
            14'd 6049: out = 12'h657;
            14'd 6050: out = 12'h657;
            14'd 6051: out = 12'h658;
            14'd 6052: out = 12'h658;
            14'd 6053: out = 12'h658;
            14'd 6054: out = 12'h658;
            14'd 6055: out = 12'h658;
            14'd 6056: out = 12'h658;
            14'd 6057: out = 12'h659;
            14'd 6058: out = 12'h659;
            14'd 6059: out = 12'h659;
            14'd 6060: out = 12'h659;
            14'd 6061: out = 12'h659;
            14'd 6062: out = 12'h659;
            14'd 6063: out = 12'h65A;
            14'd 6064: out = 12'h65A;
            14'd 6065: out = 12'h65A;
            14'd 6066: out = 12'h65A;
            14'd 6067: out = 12'h65A;
            14'd 6068: out = 12'h65A;
            14'd 6069: out = 12'h65A;
            14'd 6070: out = 12'h65B;
            14'd 6071: out = 12'h65B;
            14'd 6072: out = 12'h65B;
            14'd 6073: out = 12'h65B;
            14'd 6074: out = 12'h65B;
            14'd 6075: out = 12'h65B;
            14'd 6076: out = 12'h65C;
            14'd 6077: out = 12'h65C;
            14'd 6078: out = 12'h65C;
            14'd 6079: out = 12'h65C;
            14'd 6080: out = 12'h65C;
            14'd 6081: out = 12'h65C;
            14'd 6082: out = 12'h65D;
            14'd 6083: out = 12'h65D;
            14'd 6084: out = 12'h65D;
            14'd 6085: out = 12'h65D;
            14'd 6086: out = 12'h65D;
            14'd 6087: out = 12'h65D;
            14'd 6088: out = 12'h65D;
            14'd 6089: out = 12'h65E;
            14'd 6090: out = 12'h65E;
            14'd 6091: out = 12'h65E;
            14'd 6092: out = 12'h65E;
            14'd 6093: out = 12'h65E;
            14'd 6094: out = 12'h65E;
            14'd 6095: out = 12'h65F;
            14'd 6096: out = 12'h65F;
            14'd 6097: out = 12'h65F;
            14'd 6098: out = 12'h65F;
            14'd 6099: out = 12'h65F;
            14'd 6100: out = 12'h65F;
            14'd 6101: out = 12'h660;
            14'd 6102: out = 12'h660;
            14'd 6103: out = 12'h660;
            14'd 6104: out = 12'h660;
            14'd 6105: out = 12'h660;
            14'd 6106: out = 12'h660;
            14'd 6107: out = 12'h661;
            14'd 6108: out = 12'h661;
            14'd 6109: out = 12'h661;
            14'd 6110: out = 12'h661;
            14'd 6111: out = 12'h661;
            14'd 6112: out = 12'h661;
            14'd 6113: out = 12'h661;
            14'd 6114: out = 12'h662;
            14'd 6115: out = 12'h662;
            14'd 6116: out = 12'h662;
            14'd 6117: out = 12'h662;
            14'd 6118: out = 12'h662;
            14'd 6119: out = 12'h662;
            14'd 6120: out = 12'h663;
            14'd 6121: out = 12'h663;
            14'd 6122: out = 12'h663;
            14'd 6123: out = 12'h663;
            14'd 6124: out = 12'h663;
            14'd 6125: out = 12'h663;
            14'd 6126: out = 12'h664;
            14'd 6127: out = 12'h664;
            14'd 6128: out = 12'h664;
            14'd 6129: out = 12'h664;
            14'd 6130: out = 12'h664;
            14'd 6131: out = 12'h664;
            14'd 6132: out = 12'h664;
            14'd 6133: out = 12'h665;
            14'd 6134: out = 12'h665;
            14'd 6135: out = 12'h665;
            14'd 6136: out = 12'h665;
            14'd 6137: out = 12'h665;
            14'd 6138: out = 12'h665;
            14'd 6139: out = 12'h666;
            14'd 6140: out = 12'h666;
            14'd 6141: out = 12'h666;
            14'd 6142: out = 12'h666;
            14'd 6143: out = 12'h666;
            14'd 6144: out = 12'h666;
            14'd 6145: out = 12'h667;
            14'd 6146: out = 12'h667;
            14'd 6147: out = 12'h667;
            14'd 6148: out = 12'h667;
            14'd 6149: out = 12'h667;
            14'd 6150: out = 12'h667;
            14'd 6151: out = 12'h668;
            14'd 6152: out = 12'h668;
            14'd 6153: out = 12'h668;
            14'd 6154: out = 12'h668;
            14'd 6155: out = 12'h668;
            14'd 6156: out = 12'h668;
            14'd 6157: out = 12'h668;
            14'd 6158: out = 12'h669;
            14'd 6159: out = 12'h669;
            14'd 6160: out = 12'h669;
            14'd 6161: out = 12'h669;
            14'd 6162: out = 12'h669;
            14'd 6163: out = 12'h669;
            14'd 6164: out = 12'h66A;
            14'd 6165: out = 12'h66A;
            14'd 6166: out = 12'h66A;
            14'd 6167: out = 12'h66A;
            14'd 6168: out = 12'h66A;
            14'd 6169: out = 12'h66A;
            14'd 6170: out = 12'h66B;
            14'd 6171: out = 12'h66B;
            14'd 6172: out = 12'h66B;
            14'd 6173: out = 12'h66B;
            14'd 6174: out = 12'h66B;
            14'd 6175: out = 12'h66B;
            14'd 6176: out = 12'h66C;
            14'd 6177: out = 12'h66C;
            14'd 6178: out = 12'h66C;
            14'd 6179: out = 12'h66C;
            14'd 6180: out = 12'h66C;
            14'd 6181: out = 12'h66C;
            14'd 6182: out = 12'h66D;
            14'd 6183: out = 12'h66D;
            14'd 6184: out = 12'h66D;
            14'd 6185: out = 12'h66D;
            14'd 6186: out = 12'h66D;
            14'd 6187: out = 12'h66D;
            14'd 6188: out = 12'h66D;
            14'd 6189: out = 12'h66E;
            14'd 6190: out = 12'h66E;
            14'd 6191: out = 12'h66E;
            14'd 6192: out = 12'h66E;
            14'd 6193: out = 12'h66E;
            14'd 6194: out = 12'h66E;
            14'd 6195: out = 12'h66F;
            14'd 6196: out = 12'h66F;
            14'd 6197: out = 12'h66F;
            14'd 6198: out = 12'h66F;
            14'd 6199: out = 12'h66F;
            14'd 6200: out = 12'h66F;
            14'd 6201: out = 12'h670;
            14'd 6202: out = 12'h670;
            14'd 6203: out = 12'h670;
            14'd 6204: out = 12'h670;
            14'd 6205: out = 12'h670;
            14'd 6206: out = 12'h670;
            14'd 6207: out = 12'h671;
            14'd 6208: out = 12'h671;
            14'd 6209: out = 12'h671;
            14'd 6210: out = 12'h671;
            14'd 6211: out = 12'h671;
            14'd 6212: out = 12'h671;
            14'd 6213: out = 12'h672;
            14'd 6214: out = 12'h672;
            14'd 6215: out = 12'h672;
            14'd 6216: out = 12'h672;
            14'd 6217: out = 12'h672;
            14'd 6218: out = 12'h672;
            14'd 6219: out = 12'h672;
            14'd 6220: out = 12'h673;
            14'd 6221: out = 12'h673;
            14'd 6222: out = 12'h673;
            14'd 6223: out = 12'h673;
            14'd 6224: out = 12'h673;
            14'd 6225: out = 12'h673;
            14'd 6226: out = 12'h674;
            14'd 6227: out = 12'h674;
            14'd 6228: out = 12'h674;
            14'd 6229: out = 12'h674;
            14'd 6230: out = 12'h674;
            14'd 6231: out = 12'h674;
            14'd 6232: out = 12'h675;
            14'd 6233: out = 12'h675;
            14'd 6234: out = 12'h675;
            14'd 6235: out = 12'h675;
            14'd 6236: out = 12'h675;
            14'd 6237: out = 12'h675;
            14'd 6238: out = 12'h676;
            14'd 6239: out = 12'h676;
            14'd 6240: out = 12'h676;
            14'd 6241: out = 12'h676;
            14'd 6242: out = 12'h676;
            14'd 6243: out = 12'h676;
            14'd 6244: out = 12'h677;
            14'd 6245: out = 12'h677;
            14'd 6246: out = 12'h677;
            14'd 6247: out = 12'h677;
            14'd 6248: out = 12'h677;
            14'd 6249: out = 12'h677;
            14'd 6250: out = 12'h678;
            14'd 6251: out = 12'h678;
            14'd 6252: out = 12'h678;
            14'd 6253: out = 12'h678;
            14'd 6254: out = 12'h678;
            14'd 6255: out = 12'h678;
            14'd 6256: out = 12'h679;
            14'd 6257: out = 12'h679;
            14'd 6258: out = 12'h679;
            14'd 6259: out = 12'h679;
            14'd 6260: out = 12'h679;
            14'd 6261: out = 12'h679;
            14'd 6262: out = 12'h67A;
            14'd 6263: out = 12'h67A;
            14'd 6264: out = 12'h67A;
            14'd 6265: out = 12'h67A;
            14'd 6266: out = 12'h67A;
            14'd 6267: out = 12'h67A;
            14'd 6268: out = 12'h67A;
            14'd 6269: out = 12'h67B;
            14'd 6270: out = 12'h67B;
            14'd 6271: out = 12'h67B;
            14'd 6272: out = 12'h67B;
            14'd 6273: out = 12'h67B;
            14'd 6274: out = 12'h67B;
            14'd 6275: out = 12'h67C;
            14'd 6276: out = 12'h67C;
            14'd 6277: out = 12'h67C;
            14'd 6278: out = 12'h67C;
            14'd 6279: out = 12'h67C;
            14'd 6280: out = 12'h67C;
            14'd 6281: out = 12'h67D;
            14'd 6282: out = 12'h67D;
            14'd 6283: out = 12'h67D;
            14'd 6284: out = 12'h67D;
            14'd 6285: out = 12'h67D;
            14'd 6286: out = 12'h67D;
            14'd 6287: out = 12'h67E;
            14'd 6288: out = 12'h67E;
            14'd 6289: out = 12'h67E;
            14'd 6290: out = 12'h67E;
            14'd 6291: out = 12'h67E;
            14'd 6292: out = 12'h67E;
            14'd 6293: out = 12'h67F;
            14'd 6294: out = 12'h67F;
            14'd 6295: out = 12'h67F;
            14'd 6296: out = 12'h67F;
            14'd 6297: out = 12'h67F;
            14'd 6298: out = 12'h67F;
            14'd 6299: out = 12'h680;
            14'd 6300: out = 12'h680;
            14'd 6301: out = 12'h680;
            14'd 6302: out = 12'h680;
            14'd 6303: out = 12'h680;
            14'd 6304: out = 12'h680;
            14'd 6305: out = 12'h681;
            14'd 6306: out = 12'h681;
            14'd 6307: out = 12'h681;
            14'd 6308: out = 12'h681;
            14'd 6309: out = 12'h681;
            14'd 6310: out = 12'h681;
            14'd 6311: out = 12'h682;
            14'd 6312: out = 12'h682;
            14'd 6313: out = 12'h682;
            14'd 6314: out = 12'h682;
            14'd 6315: out = 12'h682;
            14'd 6316: out = 12'h682;
            14'd 6317: out = 12'h683;
            14'd 6318: out = 12'h683;
            14'd 6319: out = 12'h683;
            14'd 6320: out = 12'h683;
            14'd 6321: out = 12'h683;
            14'd 6322: out = 12'h683;
            14'd 6323: out = 12'h684;
            14'd 6324: out = 12'h684;
            14'd 6325: out = 12'h684;
            14'd 6326: out = 12'h684;
            14'd 6327: out = 12'h684;
            14'd 6328: out = 12'h684;
            14'd 6329: out = 12'h685;
            14'd 6330: out = 12'h685;
            14'd 6331: out = 12'h685;
            14'd 6332: out = 12'h685;
            14'd 6333: out = 12'h685;
            14'd 6334: out = 12'h685;
            14'd 6335: out = 12'h686;
            14'd 6336: out = 12'h686;
            14'd 6337: out = 12'h686;
            14'd 6338: out = 12'h686;
            14'd 6339: out = 12'h686;
            14'd 6340: out = 12'h686;
            14'd 6341: out = 12'h687;
            14'd 6342: out = 12'h687;
            14'd 6343: out = 12'h687;
            14'd 6344: out = 12'h687;
            14'd 6345: out = 12'h687;
            14'd 6346: out = 12'h687;
            14'd 6347: out = 12'h688;
            14'd 6348: out = 12'h688;
            14'd 6349: out = 12'h688;
            14'd 6350: out = 12'h688;
            14'd 6351: out = 12'h688;
            14'd 6352: out = 12'h688;
            14'd 6353: out = 12'h689;
            14'd 6354: out = 12'h689;
            14'd 6355: out = 12'h689;
            14'd 6356: out = 12'h689;
            14'd 6357: out = 12'h689;
            14'd 6358: out = 12'h689;
            14'd 6359: out = 12'h68A;
            14'd 6360: out = 12'h68A;
            14'd 6361: out = 12'h68A;
            14'd 6362: out = 12'h68A;
            14'd 6363: out = 12'h68A;
            14'd 6364: out = 12'h68A;
            14'd 6365: out = 12'h68B;
            14'd 6366: out = 12'h68B;
            14'd 6367: out = 12'h68B;
            14'd 6368: out = 12'h68B;
            14'd 6369: out = 12'h68B;
            14'd 6370: out = 12'h68B;
            14'd 6371: out = 12'h68C;
            14'd 6372: out = 12'h68C;
            14'd 6373: out = 12'h68C;
            14'd 6374: out = 12'h68C;
            14'd 6375: out = 12'h68C;
            14'd 6376: out = 12'h68C;
            14'd 6377: out = 12'h68D;
            14'd 6378: out = 12'h68D;
            14'd 6379: out = 12'h68D;
            14'd 6380: out = 12'h68D;
            14'd 6381: out = 12'h68D;
            14'd 6382: out = 12'h68D;
            14'd 6383: out = 12'h68E;
            14'd 6384: out = 12'h68E;
            14'd 6385: out = 12'h68E;
            14'd 6386: out = 12'h68E;
            14'd 6387: out = 12'h68E;
            14'd 6388: out = 12'h68E;
            14'd 6389: out = 12'h68F;
            14'd 6390: out = 12'h68F;
            14'd 6391: out = 12'h68F;
            14'd 6392: out = 12'h68F;
            14'd 6393: out = 12'h68F;
            14'd 6394: out = 12'h68F;
            14'd 6395: out = 12'h690;
            14'd 6396: out = 12'h690;
            14'd 6397: out = 12'h690;
            14'd 6398: out = 12'h690;
            14'd 6399: out = 12'h690;
            14'd 6400: out = 12'h690;
            14'd 6401: out = 12'h691;
            14'd 6402: out = 12'h691;
            14'd 6403: out = 12'h691;
            14'd 6404: out = 12'h691;
            14'd 6405: out = 12'h691;
            14'd 6406: out = 12'h691;
            14'd 6407: out = 12'h692;
            14'd 6408: out = 12'h692;
            14'd 6409: out = 12'h692;
            14'd 6410: out = 12'h692;
            14'd 6411: out = 12'h692;
            14'd 6412: out = 12'h692;
            14'd 6413: out = 12'h693;
            14'd 6414: out = 12'h693;
            14'd 6415: out = 12'h693;
            14'd 6416: out = 12'h693;
            14'd 6417: out = 12'h693;
            14'd 6418: out = 12'h693;
            14'd 6419: out = 12'h694;
            14'd 6420: out = 12'h694;
            14'd 6421: out = 12'h694;
            14'd 6422: out = 12'h694;
            14'd 6423: out = 12'h694;
            14'd 6424: out = 12'h694;
            14'd 6425: out = 12'h695;
            14'd 6426: out = 12'h695;
            14'd 6427: out = 12'h695;
            14'd 6428: out = 12'h695;
            14'd 6429: out = 12'h695;
            14'd 6430: out = 12'h695;
            14'd 6431: out = 12'h696;
            14'd 6432: out = 12'h696;
            14'd 6433: out = 12'h696;
            14'd 6434: out = 12'h696;
            14'd 6435: out = 12'h696;
            14'd 6436: out = 12'h696;
            14'd 6437: out = 12'h697;
            14'd 6438: out = 12'h697;
            14'd 6439: out = 12'h697;
            14'd 6440: out = 12'h697;
            14'd 6441: out = 12'h697;
            14'd 6442: out = 12'h698;
            14'd 6443: out = 12'h698;
            14'd 6444: out = 12'h698;
            14'd 6445: out = 12'h698;
            14'd 6446: out = 12'h698;
            14'd 6447: out = 12'h698;
            14'd 6448: out = 12'h699;
            14'd 6449: out = 12'h699;
            14'd 6450: out = 12'h699;
            14'd 6451: out = 12'h699;
            14'd 6452: out = 12'h699;
            14'd 6453: out = 12'h699;
            14'd 6454: out = 12'h69A;
            14'd 6455: out = 12'h69A;
            14'd 6456: out = 12'h69A;
            14'd 6457: out = 12'h69A;
            14'd 6458: out = 12'h69A;
            14'd 6459: out = 12'h69A;
            14'd 6460: out = 12'h69B;
            14'd 6461: out = 12'h69B;
            14'd 6462: out = 12'h69B;
            14'd 6463: out = 12'h69B;
            14'd 6464: out = 12'h69B;
            14'd 6465: out = 12'h69B;
            14'd 6466: out = 12'h69C;
            14'd 6467: out = 12'h69C;
            14'd 6468: out = 12'h69C;
            14'd 6469: out = 12'h69C;
            14'd 6470: out = 12'h69C;
            14'd 6471: out = 12'h69C;
            14'd 6472: out = 12'h69D;
            14'd 6473: out = 12'h69D;
            14'd 6474: out = 12'h69D;
            14'd 6475: out = 12'h69D;
            14'd 6476: out = 12'h69D;
            14'd 6477: out = 12'h69D;
            14'd 6478: out = 12'h69E;
            14'd 6479: out = 12'h69E;
            14'd 6480: out = 12'h69E;
            14'd 6481: out = 12'h69E;
            14'd 6482: out = 12'h69E;
            14'd 6483: out = 12'h69E;
            14'd 6484: out = 12'h69F;
            14'd 6485: out = 12'h69F;
            14'd 6486: out = 12'h69F;
            14'd 6487: out = 12'h69F;
            14'd 6488: out = 12'h69F;
            14'd 6489: out = 12'h6A0;
            14'd 6490: out = 12'h6A0;
            14'd 6491: out = 12'h6A0;
            14'd 6492: out = 12'h6A0;
            14'd 6493: out = 12'h6A0;
            14'd 6494: out = 12'h6A0;
            14'd 6495: out = 12'h6A1;
            14'd 6496: out = 12'h6A1;
            14'd 6497: out = 12'h6A1;
            14'd 6498: out = 12'h6A1;
            14'd 6499: out = 12'h6A1;
            14'd 6500: out = 12'h6A1;
            14'd 6501: out = 12'h6A2;
            14'd 6502: out = 12'h6A2;
            14'd 6503: out = 12'h6A2;
            14'd 6504: out = 12'h6A2;
            14'd 6505: out = 12'h6A2;
            14'd 6506: out = 12'h6A2;
            14'd 6507: out = 12'h6A3;
            14'd 6508: out = 12'h6A3;
            14'd 6509: out = 12'h6A3;
            14'd 6510: out = 12'h6A3;
            14'd 6511: out = 12'h6A3;
            14'd 6512: out = 12'h6A3;
            14'd 6513: out = 12'h6A4;
            14'd 6514: out = 12'h6A4;
            14'd 6515: out = 12'h6A4;
            14'd 6516: out = 12'h6A4;
            14'd 6517: out = 12'h6A4;
            14'd 6518: out = 12'h6A5;
            14'd 6519: out = 12'h6A5;
            14'd 6520: out = 12'h6A5;
            14'd 6521: out = 12'h6A5;
            14'd 6522: out = 12'h6A5;
            14'd 6523: out = 12'h6A5;
            14'd 6524: out = 12'h6A6;
            14'd 6525: out = 12'h6A6;
            14'd 6526: out = 12'h6A6;
            14'd 6527: out = 12'h6A6;
            14'd 6528: out = 12'h6A6;
            14'd 6529: out = 12'h6A6;
            14'd 6530: out = 12'h6A7;
            14'd 6531: out = 12'h6A7;
            14'd 6532: out = 12'h6A7;
            14'd 6533: out = 12'h6A7;
            14'd 6534: out = 12'h6A7;
            14'd 6535: out = 12'h6A7;
            14'd 6536: out = 12'h6A8;
            14'd 6537: out = 12'h6A8;
            14'd 6538: out = 12'h6A8;
            14'd 6539: out = 12'h6A8;
            14'd 6540: out = 12'h6A8;
            14'd 6541: out = 12'h6A8;
            14'd 6542: out = 12'h6A9;
            14'd 6543: out = 12'h6A9;
            14'd 6544: out = 12'h6A9;
            14'd 6545: out = 12'h6A9;
            14'd 6546: out = 12'h6A9;
            14'd 6547: out = 12'h6AA;
            14'd 6548: out = 12'h6AA;
            14'd 6549: out = 12'h6AA;
            14'd 6550: out = 12'h6AA;
            14'd 6551: out = 12'h6AA;
            14'd 6552: out = 12'h6AA;
            14'd 6553: out = 12'h6AB;
            14'd 6554: out = 12'h6AB;
            14'd 6555: out = 12'h6AB;
            14'd 6556: out = 12'h6AB;
            14'd 6557: out = 12'h6AB;
            14'd 6558: out = 12'h6AB;
            14'd 6559: out = 12'h6AC;
            14'd 6560: out = 12'h6AC;
            14'd 6561: out = 12'h6AC;
            14'd 6562: out = 12'h6AC;
            14'd 6563: out = 12'h6AC;
            14'd 6564: out = 12'h6AC;
            14'd 6565: out = 12'h6AD;
            14'd 6566: out = 12'h6AD;
            14'd 6567: out = 12'h6AD;
            14'd 6568: out = 12'h6AD;
            14'd 6569: out = 12'h6AD;
            14'd 6570: out = 12'h6AE;
            14'd 6571: out = 12'h6AE;
            14'd 6572: out = 12'h6AE;
            14'd 6573: out = 12'h6AE;
            14'd 6574: out = 12'h6AE;
            14'd 6575: out = 12'h6AE;
            14'd 6576: out = 12'h6AF;
            14'd 6577: out = 12'h6AF;
            14'd 6578: out = 12'h6AF;
            14'd 6579: out = 12'h6AF;
            14'd 6580: out = 12'h6AF;
            14'd 6581: out = 12'h6AF;
            14'd 6582: out = 12'h6B0;
            14'd 6583: out = 12'h6B0;
            14'd 6584: out = 12'h6B0;
            14'd 6585: out = 12'h6B0;
            14'd 6586: out = 12'h6B0;
            14'd 6587: out = 12'h6B0;
            14'd 6588: out = 12'h6B1;
            14'd 6589: out = 12'h6B1;
            14'd 6590: out = 12'h6B1;
            14'd 6591: out = 12'h6B1;
            14'd 6592: out = 12'h6B1;
            14'd 6593: out = 12'h6B2;
            14'd 6594: out = 12'h6B2;
            14'd 6595: out = 12'h6B2;
            14'd 6596: out = 12'h6B2;
            14'd 6597: out = 12'h6B2;
            14'd 6598: out = 12'h6B2;
            14'd 6599: out = 12'h6B3;
            14'd 6600: out = 12'h6B3;
            14'd 6601: out = 12'h6B3;
            14'd 6602: out = 12'h6B3;
            14'd 6603: out = 12'h6B3;
            14'd 6604: out = 12'h6B3;
            14'd 6605: out = 12'h6B4;
            14'd 6606: out = 12'h6B4;
            14'd 6607: out = 12'h6B4;
            14'd 6608: out = 12'h6B4;
            14'd 6609: out = 12'h6B4;
            14'd 6610: out = 12'h6B5;
            14'd 6611: out = 12'h6B5;
            14'd 6612: out = 12'h6B5;
            14'd 6613: out = 12'h6B5;
            14'd 6614: out = 12'h6B5;
            14'd 6615: out = 12'h6B5;
            14'd 6616: out = 12'h6B6;
            14'd 6617: out = 12'h6B6;
            14'd 6618: out = 12'h6B6;
            14'd 6619: out = 12'h6B6;
            14'd 6620: out = 12'h6B6;
            14'd 6621: out = 12'h6B6;
            14'd 6622: out = 12'h6B7;
            14'd 6623: out = 12'h6B7;
            14'd 6624: out = 12'h6B7;
            14'd 6625: out = 12'h6B7;
            14'd 6626: out = 12'h6B7;
            14'd 6627: out = 12'h6B8;
            14'd 6628: out = 12'h6B8;
            14'd 6629: out = 12'h6B8;
            14'd 6630: out = 12'h6B8;
            14'd 6631: out = 12'h6B8;
            14'd 6632: out = 12'h6B8;
            14'd 6633: out = 12'h6B9;
            14'd 6634: out = 12'h6B9;
            14'd 6635: out = 12'h6B9;
            14'd 6636: out = 12'h6B9;
            14'd 6637: out = 12'h6B9;
            14'd 6638: out = 12'h6B9;
            14'd 6639: out = 12'h6BA;
            14'd 6640: out = 12'h6BA;
            14'd 6641: out = 12'h6BA;
            14'd 6642: out = 12'h6BA;
            14'd 6643: out = 12'h6BA;
            14'd 6644: out = 12'h6BB;
            14'd 6645: out = 12'h6BB;
            14'd 6646: out = 12'h6BB;
            14'd 6647: out = 12'h6BB;
            14'd 6648: out = 12'h6BB;
            14'd 6649: out = 12'h6BB;
            14'd 6650: out = 12'h6BC;
            14'd 6651: out = 12'h6BC;
            14'd 6652: out = 12'h6BC;
            14'd 6653: out = 12'h6BC;
            14'd 6654: out = 12'h6BC;
            14'd 6655: out = 12'h6BC;
            14'd 6656: out = 12'h6BD;
            14'd 6657: out = 12'h6BD;
            14'd 6658: out = 12'h6BD;
            14'd 6659: out = 12'h6BD;
            14'd 6660: out = 12'h6BD;
            14'd 6661: out = 12'h6BE;
            14'd 6662: out = 12'h6BE;
            14'd 6663: out = 12'h6BE;
            14'd 6664: out = 12'h6BE;
            14'd 6665: out = 12'h6BE;
            14'd 6666: out = 12'h6BE;
            14'd 6667: out = 12'h6BF;
            14'd 6668: out = 12'h6BF;
            14'd 6669: out = 12'h6BF;
            14'd 6670: out = 12'h6BF;
            14'd 6671: out = 12'h6BF;
            14'd 6672: out = 12'h6BF;
            14'd 6673: out = 12'h6C0;
            14'd 6674: out = 12'h6C0;
            14'd 6675: out = 12'h6C0;
            14'd 6676: out = 12'h6C0;
            14'd 6677: out = 12'h6C0;
            14'd 6678: out = 12'h6C1;
            14'd 6679: out = 12'h6C1;
            14'd 6680: out = 12'h6C1;
            14'd 6681: out = 12'h6C1;
            14'd 6682: out = 12'h6C1;
            14'd 6683: out = 12'h6C1;
            14'd 6684: out = 12'h6C2;
            14'd 6685: out = 12'h6C2;
            14'd 6686: out = 12'h6C2;
            14'd 6687: out = 12'h6C2;
            14'd 6688: out = 12'h6C2;
            14'd 6689: out = 12'h6C3;
            14'd 6690: out = 12'h6C3;
            14'd 6691: out = 12'h6C3;
            14'd 6692: out = 12'h6C3;
            14'd 6693: out = 12'h6C3;
            14'd 6694: out = 12'h6C3;
            14'd 6695: out = 12'h6C4;
            14'd 6696: out = 12'h6C4;
            14'd 6697: out = 12'h6C4;
            14'd 6698: out = 12'h6C4;
            14'd 6699: out = 12'h6C4;
            14'd 6700: out = 12'h6C4;
            14'd 6701: out = 12'h6C5;
            14'd 6702: out = 12'h6C5;
            14'd 6703: out = 12'h6C5;
            14'd 6704: out = 12'h6C5;
            14'd 6705: out = 12'h6C5;
            14'd 6706: out = 12'h6C6;
            14'd 6707: out = 12'h6C6;
            14'd 6708: out = 12'h6C6;
            14'd 6709: out = 12'h6C6;
            14'd 6710: out = 12'h6C6;
            14'd 6711: out = 12'h6C6;
            14'd 6712: out = 12'h6C7;
            14'd 6713: out = 12'h6C7;
            14'd 6714: out = 12'h6C7;
            14'd 6715: out = 12'h6C7;
            14'd 6716: out = 12'h6C7;
            14'd 6717: out = 12'h6C8;
            14'd 6718: out = 12'h6C8;
            14'd 6719: out = 12'h6C8;
            14'd 6720: out = 12'h6C8;
            14'd 6721: out = 12'h6C8;
            14'd 6722: out = 12'h6C8;
            14'd 6723: out = 12'h6C9;
            14'd 6724: out = 12'h6C9;
            14'd 6725: out = 12'h6C9;
            14'd 6726: out = 12'h6C9;
            14'd 6727: out = 12'h6C9;
            14'd 6728: out = 12'h6C9;
            14'd 6729: out = 12'h6CA;
            14'd 6730: out = 12'h6CA;
            14'd 6731: out = 12'h6CA;
            14'd 6732: out = 12'h6CA;
            14'd 6733: out = 12'h6CA;
            14'd 6734: out = 12'h6CB;
            14'd 6735: out = 12'h6CB;
            14'd 6736: out = 12'h6CB;
            14'd 6737: out = 12'h6CB;
            14'd 6738: out = 12'h6CB;
            14'd 6739: out = 12'h6CB;
            14'd 6740: out = 12'h6CC;
            14'd 6741: out = 12'h6CC;
            14'd 6742: out = 12'h6CC;
            14'd 6743: out = 12'h6CC;
            14'd 6744: out = 12'h6CC;
            14'd 6745: out = 12'h6CD;
            14'd 6746: out = 12'h6CD;
            14'd 6747: out = 12'h6CD;
            14'd 6748: out = 12'h6CD;
            14'd 6749: out = 12'h6CD;
            14'd 6750: out = 12'h6CD;
            14'd 6751: out = 12'h6CE;
            14'd 6752: out = 12'h6CE;
            14'd 6753: out = 12'h6CE;
            14'd 6754: out = 12'h6CE;
            14'd 6755: out = 12'h6CE;
            14'd 6756: out = 12'h6CF;
            14'd 6757: out = 12'h6CF;
            14'd 6758: out = 12'h6CF;
            14'd 6759: out = 12'h6CF;
            14'd 6760: out = 12'h6CF;
            14'd 6761: out = 12'h6CF;
            14'd 6762: out = 12'h6D0;
            14'd 6763: out = 12'h6D0;
            14'd 6764: out = 12'h6D0;
            14'd 6765: out = 12'h6D0;
            14'd 6766: out = 12'h6D0;
            14'd 6767: out = 12'h6D1;
            14'd 6768: out = 12'h6D1;
            14'd 6769: out = 12'h6D1;
            14'd 6770: out = 12'h6D1;
            14'd 6771: out = 12'h6D1;
            14'd 6772: out = 12'h6D1;
            14'd 6773: out = 12'h6D2;
            14'd 6774: out = 12'h6D2;
            14'd 6775: out = 12'h6D2;
            14'd 6776: out = 12'h6D2;
            14'd 6777: out = 12'h6D2;
            14'd 6778: out = 12'h6D3;
            14'd 6779: out = 12'h6D3;
            14'd 6780: out = 12'h6D3;
            14'd 6781: out = 12'h6D3;
            14'd 6782: out = 12'h6D3;
            14'd 6783: out = 12'h6D3;
            14'd 6784: out = 12'h6D4;
            14'd 6785: out = 12'h6D4;
            14'd 6786: out = 12'h6D4;
            14'd 6787: out = 12'h6D4;
            14'd 6788: out = 12'h6D4;
            14'd 6789: out = 12'h6D5;
            14'd 6790: out = 12'h6D5;
            14'd 6791: out = 12'h6D5;
            14'd 6792: out = 12'h6D5;
            14'd 6793: out = 12'h6D5;
            14'd 6794: out = 12'h6D5;
            14'd 6795: out = 12'h6D6;
            14'd 6796: out = 12'h6D6;
            14'd 6797: out = 12'h6D6;
            14'd 6798: out = 12'h6D6;
            14'd 6799: out = 12'h6D6;
            14'd 6800: out = 12'h6D7;
            14'd 6801: out = 12'h6D7;
            14'd 6802: out = 12'h6D7;
            14'd 6803: out = 12'h6D7;
            14'd 6804: out = 12'h6D7;
            14'd 6805: out = 12'h6D7;
            14'd 6806: out = 12'h6D8;
            14'd 6807: out = 12'h6D8;
            14'd 6808: out = 12'h6D8;
            14'd 6809: out = 12'h6D8;
            14'd 6810: out = 12'h6D8;
            14'd 6811: out = 12'h6D9;
            14'd 6812: out = 12'h6D9;
            14'd 6813: out = 12'h6D9;
            14'd 6814: out = 12'h6D9;
            14'd 6815: out = 12'h6D9;
            14'd 6816: out = 12'h6D9;
            14'd 6817: out = 12'h6DA;
            14'd 6818: out = 12'h6DA;
            14'd 6819: out = 12'h6DA;
            14'd 6820: out = 12'h6DA;
            14'd 6821: out = 12'h6DA;
            14'd 6822: out = 12'h6DB;
            14'd 6823: out = 12'h6DB;
            14'd 6824: out = 12'h6DB;
            14'd 6825: out = 12'h6DB;
            14'd 6826: out = 12'h6DB;
            14'd 6827: out = 12'h6DB;
            14'd 6828: out = 12'h6DC;
            14'd 6829: out = 12'h6DC;
            14'd 6830: out = 12'h6DC;
            14'd 6831: out = 12'h6DC;
            14'd 6832: out = 12'h6DC;
            14'd 6833: out = 12'h6DD;
            14'd 6834: out = 12'h6DD;
            14'd 6835: out = 12'h6DD;
            14'd 6836: out = 12'h6DD;
            14'd 6837: out = 12'h6DD;
            14'd 6838: out = 12'h6DE;
            14'd 6839: out = 12'h6DE;
            14'd 6840: out = 12'h6DE;
            14'd 6841: out = 12'h6DE;
            14'd 6842: out = 12'h6DE;
            14'd 6843: out = 12'h6DE;
            14'd 6844: out = 12'h6DF;
            14'd 6845: out = 12'h6DF;
            14'd 6846: out = 12'h6DF;
            14'd 6847: out = 12'h6DF;
            14'd 6848: out = 12'h6DF;
            14'd 6849: out = 12'h6E0;
            14'd 6850: out = 12'h6E0;
            14'd 6851: out = 12'h6E0;
            14'd 6852: out = 12'h6E0;
            14'd 6853: out = 12'h6E0;
            14'd 6854: out = 12'h6E0;
            14'd 6855: out = 12'h6E1;
            14'd 6856: out = 12'h6E1;
            14'd 6857: out = 12'h6E1;
            14'd 6858: out = 12'h6E1;
            14'd 6859: out = 12'h6E1;
            14'd 6860: out = 12'h6E2;
            14'd 6861: out = 12'h6E2;
            14'd 6862: out = 12'h6E2;
            14'd 6863: out = 12'h6E2;
            14'd 6864: out = 12'h6E2;
            14'd 6865: out = 12'h6E2;
            14'd 6866: out = 12'h6E3;
            14'd 6867: out = 12'h6E3;
            14'd 6868: out = 12'h6E3;
            14'd 6869: out = 12'h6E3;
            14'd 6870: out = 12'h6E3;
            14'd 6871: out = 12'h6E4;
            14'd 6872: out = 12'h6E4;
            14'd 6873: out = 12'h6E4;
            14'd 6874: out = 12'h6E4;
            14'd 6875: out = 12'h6E4;
            14'd 6876: out = 12'h6E5;
            14'd 6877: out = 12'h6E5;
            14'd 6878: out = 12'h6E5;
            14'd 6879: out = 12'h6E5;
            14'd 6880: out = 12'h6E5;
            14'd 6881: out = 12'h6E5;
            14'd 6882: out = 12'h6E6;
            14'd 6883: out = 12'h6E6;
            14'd 6884: out = 12'h6E6;
            14'd 6885: out = 12'h6E6;
            14'd 6886: out = 12'h6E6;
            14'd 6887: out = 12'h6E7;
            14'd 6888: out = 12'h6E7;
            14'd 6889: out = 12'h6E7;
            14'd 6890: out = 12'h6E7;
            14'd 6891: out = 12'h6E7;
            14'd 6892: out = 12'h6E8;
            14'd 6893: out = 12'h6E8;
            14'd 6894: out = 12'h6E8;
            14'd 6895: out = 12'h6E8;
            14'd 6896: out = 12'h6E8;
            14'd 6897: out = 12'h6E8;
            14'd 6898: out = 12'h6E9;
            14'd 6899: out = 12'h6E9;
            14'd 6900: out = 12'h6E9;
            14'd 6901: out = 12'h6E9;
            14'd 6902: out = 12'h6E9;
            14'd 6903: out = 12'h6EA;
            14'd 6904: out = 12'h6EA;
            14'd 6905: out = 12'h6EA;
            14'd 6906: out = 12'h6EA;
            14'd 6907: out = 12'h6EA;
            14'd 6908: out = 12'h6EA;
            14'd 6909: out = 12'h6EB;
            14'd 6910: out = 12'h6EB;
            14'd 6911: out = 12'h6EB;
            14'd 6912: out = 12'h6EB;
            14'd 6913: out = 12'h6EB;
            14'd 6914: out = 12'h6EC;
            14'd 6915: out = 12'h6EC;
            14'd 6916: out = 12'h6EC;
            14'd 6917: out = 12'h6EC;
            14'd 6918: out = 12'h6EC;
            14'd 6919: out = 12'h6ED;
            14'd 6920: out = 12'h6ED;
            14'd 6921: out = 12'h6ED;
            14'd 6922: out = 12'h6ED;
            14'd 6923: out = 12'h6ED;
            14'd 6924: out = 12'h6ED;
            14'd 6925: out = 12'h6EE;
            14'd 6926: out = 12'h6EE;
            14'd 6927: out = 12'h6EE;
            14'd 6928: out = 12'h6EE;
            14'd 6929: out = 12'h6EE;
            14'd 6930: out = 12'h6EF;
            14'd 6931: out = 12'h6EF;
            14'd 6932: out = 12'h6EF;
            14'd 6933: out = 12'h6EF;
            14'd 6934: out = 12'h6EF;
            14'd 6935: out = 12'h6F0;
            14'd 6936: out = 12'h6F0;
            14'd 6937: out = 12'h6F0;
            14'd 6938: out = 12'h6F0;
            14'd 6939: out = 12'h6F0;
            14'd 6940: out = 12'h6F0;
            14'd 6941: out = 12'h6F1;
            14'd 6942: out = 12'h6F1;
            14'd 6943: out = 12'h6F1;
            14'd 6944: out = 12'h6F1;
            14'd 6945: out = 12'h6F1;
            14'd 6946: out = 12'h6F2;
            14'd 6947: out = 12'h6F2;
            14'd 6948: out = 12'h6F2;
            14'd 6949: out = 12'h6F2;
            14'd 6950: out = 12'h6F2;
            14'd 6951: out = 12'h6F3;
            14'd 6952: out = 12'h6F3;
            14'd 6953: out = 12'h6F3;
            14'd 6954: out = 12'h6F3;
            14'd 6955: out = 12'h6F3;
            14'd 6956: out = 12'h6F4;
            14'd 6957: out = 12'h6F4;
            14'd 6958: out = 12'h6F4;
            14'd 6959: out = 12'h6F4;
            14'd 6960: out = 12'h6F4;
            14'd 6961: out = 12'h6F4;
            14'd 6962: out = 12'h6F5;
            14'd 6963: out = 12'h6F5;
            14'd 6964: out = 12'h6F5;
            14'd 6965: out = 12'h6F5;
            14'd 6966: out = 12'h6F5;
            14'd 6967: out = 12'h6F6;
            14'd 6968: out = 12'h6F6;
            14'd 6969: out = 12'h6F6;
            14'd 6970: out = 12'h6F6;
            14'd 6971: out = 12'h6F6;
            14'd 6972: out = 12'h6F7;
            14'd 6973: out = 12'h6F7;
            14'd 6974: out = 12'h6F7;
            14'd 6975: out = 12'h6F7;
            14'd 6976: out = 12'h6F7;
            14'd 6977: out = 12'h6F7;
            14'd 6978: out = 12'h6F8;
            14'd 6979: out = 12'h6F8;
            14'd 6980: out = 12'h6F8;
            14'd 6981: out = 12'h6F8;
            14'd 6982: out = 12'h6F8;
            14'd 6983: out = 12'h6F9;
            14'd 6984: out = 12'h6F9;
            14'd 6985: out = 12'h6F9;
            14'd 6986: out = 12'h6F9;
            14'd 6987: out = 12'h6F9;
            14'd 6988: out = 12'h6FA;
            14'd 6989: out = 12'h6FA;
            14'd 6990: out = 12'h6FA;
            14'd 6991: out = 12'h6FA;
            14'd 6992: out = 12'h6FA;
            14'd 6993: out = 12'h6FB;
            14'd 6994: out = 12'h6FB;
            14'd 6995: out = 12'h6FB;
            14'd 6996: out = 12'h6FB;
            14'd 6997: out = 12'h6FB;
            14'd 6998: out = 12'h6FB;
            14'd 6999: out = 12'h6FC;
            14'd 7000: out = 12'h6FC;
            14'd 7001: out = 12'h6FC;
            14'd 7002: out = 12'h6FC;
            14'd 7003: out = 12'h6FC;
            14'd 7004: out = 12'h6FD;
            14'd 7005: out = 12'h6FD;
            14'd 7006: out = 12'h6FD;
            14'd 7007: out = 12'h6FD;
            14'd 7008: out = 12'h6FD;
            14'd 7009: out = 12'h6FE;
            14'd 7010: out = 12'h6FE;
            14'd 7011: out = 12'h6FE;
            14'd 7012: out = 12'h6FE;
            14'd 7013: out = 12'h6FE;
            14'd 7014: out = 12'h6FF;
            14'd 7015: out = 12'h6FF;
            14'd 7016: out = 12'h6FF;
            14'd 7017: out = 12'h6FF;
            14'd 7018: out = 12'h6FF;
            14'd 7019: out = 12'h6FF;
            14'd 7020: out = 12'h700;
            14'd 7021: out = 12'h700;
            14'd 7022: out = 12'h700;
            14'd 7023: out = 12'h700;
            14'd 7024: out = 12'h700;
            14'd 7025: out = 12'h701;
            14'd 7026: out = 12'h701;
            14'd 7027: out = 12'h701;
            14'd 7028: out = 12'h701;
            14'd 7029: out = 12'h701;
            14'd 7030: out = 12'h702;
            14'd 7031: out = 12'h702;
            14'd 7032: out = 12'h702;
            14'd 7033: out = 12'h702;
            14'd 7034: out = 12'h702;
            14'd 7035: out = 12'h703;
            14'd 7036: out = 12'h703;
            14'd 7037: out = 12'h703;
            14'd 7038: out = 12'h703;
            14'd 7039: out = 12'h703;
            14'd 7040: out = 12'h704;
            14'd 7041: out = 12'h704;
            14'd 7042: out = 12'h704;
            14'd 7043: out = 12'h704;
            14'd 7044: out = 12'h704;
            14'd 7045: out = 12'h704;
            14'd 7046: out = 12'h705;
            14'd 7047: out = 12'h705;
            14'd 7048: out = 12'h705;
            14'd 7049: out = 12'h705;
            14'd 7050: out = 12'h705;
            14'd 7051: out = 12'h706;
            14'd 7052: out = 12'h706;
            14'd 7053: out = 12'h706;
            14'd 7054: out = 12'h706;
            14'd 7055: out = 12'h706;
            14'd 7056: out = 12'h707;
            14'd 7057: out = 12'h707;
            14'd 7058: out = 12'h707;
            14'd 7059: out = 12'h707;
            14'd 7060: out = 12'h707;
            14'd 7061: out = 12'h708;
            14'd 7062: out = 12'h708;
            14'd 7063: out = 12'h708;
            14'd 7064: out = 12'h708;
            14'd 7065: out = 12'h708;
            14'd 7066: out = 12'h709;
            14'd 7067: out = 12'h709;
            14'd 7068: out = 12'h709;
            14'd 7069: out = 12'h709;
            14'd 7070: out = 12'h709;
            14'd 7071: out = 12'h709;
            14'd 7072: out = 12'h70A;
            14'd 7073: out = 12'h70A;
            14'd 7074: out = 12'h70A;
            14'd 7075: out = 12'h70A;
            14'd 7076: out = 12'h70A;
            14'd 7077: out = 12'h70B;
            14'd 7078: out = 12'h70B;
            14'd 7079: out = 12'h70B;
            14'd 7080: out = 12'h70B;
            14'd 7081: out = 12'h70B;
            14'd 7082: out = 12'h70C;
            14'd 7083: out = 12'h70C;
            14'd 7084: out = 12'h70C;
            14'd 7085: out = 12'h70C;
            14'd 7086: out = 12'h70C;
            14'd 7087: out = 12'h70D;
            14'd 7088: out = 12'h70D;
            14'd 7089: out = 12'h70D;
            14'd 7090: out = 12'h70D;
            14'd 7091: out = 12'h70D;
            14'd 7092: out = 12'h70E;
            14'd 7093: out = 12'h70E;
            14'd 7094: out = 12'h70E;
            14'd 7095: out = 12'h70E;
            14'd 7096: out = 12'h70E;
            14'd 7097: out = 12'h70F;
            14'd 7098: out = 12'h70F;
            14'd 7099: out = 12'h70F;
            14'd 7100: out = 12'h70F;
            14'd 7101: out = 12'h70F;
            14'd 7102: out = 12'h710;
            14'd 7103: out = 12'h710;
            14'd 7104: out = 12'h710;
            14'd 7105: out = 12'h710;
            14'd 7106: out = 12'h710;
            14'd 7107: out = 12'h710;
            14'd 7108: out = 12'h711;
            14'd 7109: out = 12'h711;
            14'd 7110: out = 12'h711;
            14'd 7111: out = 12'h711;
            14'd 7112: out = 12'h711;
            14'd 7113: out = 12'h712;
            14'd 7114: out = 12'h712;
            14'd 7115: out = 12'h712;
            14'd 7116: out = 12'h712;
            14'd 7117: out = 12'h712;
            14'd 7118: out = 12'h713;
            14'd 7119: out = 12'h713;
            14'd 7120: out = 12'h713;
            14'd 7121: out = 12'h713;
            14'd 7122: out = 12'h713;
            14'd 7123: out = 12'h714;
            14'd 7124: out = 12'h714;
            14'd 7125: out = 12'h714;
            14'd 7126: out = 12'h714;
            14'd 7127: out = 12'h714;
            14'd 7128: out = 12'h715;
            14'd 7129: out = 12'h715;
            14'd 7130: out = 12'h715;
            14'd 7131: out = 12'h715;
            14'd 7132: out = 12'h715;
            14'd 7133: out = 12'h716;
            14'd 7134: out = 12'h716;
            14'd 7135: out = 12'h716;
            14'd 7136: out = 12'h716;
            14'd 7137: out = 12'h716;
            14'd 7138: out = 12'h717;
            14'd 7139: out = 12'h717;
            14'd 7140: out = 12'h717;
            14'd 7141: out = 12'h717;
            14'd 7142: out = 12'h717;
            14'd 7143: out = 12'h718;
            14'd 7144: out = 12'h718;
            14'd 7145: out = 12'h718;
            14'd 7146: out = 12'h718;
            14'd 7147: out = 12'h718;
            14'd 7148: out = 12'h719;
            14'd 7149: out = 12'h719;
            14'd 7150: out = 12'h719;
            14'd 7151: out = 12'h719;
            14'd 7152: out = 12'h719;
            14'd 7153: out = 12'h719;
            14'd 7154: out = 12'h71A;
            14'd 7155: out = 12'h71A;
            14'd 7156: out = 12'h71A;
            14'd 7157: out = 12'h71A;
            14'd 7158: out = 12'h71A;
            14'd 7159: out = 12'h71B;
            14'd 7160: out = 12'h71B;
            14'd 7161: out = 12'h71B;
            14'd 7162: out = 12'h71B;
            14'd 7163: out = 12'h71B;
            14'd 7164: out = 12'h71C;
            14'd 7165: out = 12'h71C;
            14'd 7166: out = 12'h71C;
            14'd 7167: out = 12'h71C;
            14'd 7168: out = 12'h71C;
            14'd 7169: out = 12'h71D;
            14'd 7170: out = 12'h71D;
            14'd 7171: out = 12'h71D;
            14'd 7172: out = 12'h71D;
            14'd 7173: out = 12'h71D;
            14'd 7174: out = 12'h71E;
            14'd 7175: out = 12'h71E;
            14'd 7176: out = 12'h71E;
            14'd 7177: out = 12'h71E;
            14'd 7178: out = 12'h71E;
            14'd 7179: out = 12'h71F;
            14'd 7180: out = 12'h71F;
            14'd 7181: out = 12'h71F;
            14'd 7182: out = 12'h71F;
            14'd 7183: out = 12'h71F;
            14'd 7184: out = 12'h720;
            14'd 7185: out = 12'h720;
            14'd 7186: out = 12'h720;
            14'd 7187: out = 12'h720;
            14'd 7188: out = 12'h720;
            14'd 7189: out = 12'h721;
            14'd 7190: out = 12'h721;
            14'd 7191: out = 12'h721;
            14'd 7192: out = 12'h721;
            14'd 7193: out = 12'h721;
            14'd 7194: out = 12'h722;
            14'd 7195: out = 12'h722;
            14'd 7196: out = 12'h722;
            14'd 7197: out = 12'h722;
            14'd 7198: out = 12'h722;
            14'd 7199: out = 12'h723;
            14'd 7200: out = 12'h723;
            14'd 7201: out = 12'h723;
            14'd 7202: out = 12'h723;
            14'd 7203: out = 12'h723;
            14'd 7204: out = 12'h724;
            14'd 7205: out = 12'h724;
            14'd 7206: out = 12'h724;
            14'd 7207: out = 12'h724;
            14'd 7208: out = 12'h724;
            14'd 7209: out = 12'h725;
            14'd 7210: out = 12'h725;
            14'd 7211: out = 12'h725;
            14'd 7212: out = 12'h725;
            14'd 7213: out = 12'h725;
            14'd 7214: out = 12'h726;
            14'd 7215: out = 12'h726;
            14'd 7216: out = 12'h726;
            14'd 7217: out = 12'h726;
            14'd 7218: out = 12'h726;
            14'd 7219: out = 12'h727;
            14'd 7220: out = 12'h727;
            14'd 7221: out = 12'h727;
            14'd 7222: out = 12'h727;
            14'd 7223: out = 12'h727;
            14'd 7224: out = 12'h728;
            14'd 7225: out = 12'h728;
            14'd 7226: out = 12'h728;
            14'd 7227: out = 12'h728;
            14'd 7228: out = 12'h728;
            14'd 7229: out = 12'h729;
            14'd 7230: out = 12'h729;
            14'd 7231: out = 12'h729;
            14'd 7232: out = 12'h729;
            14'd 7233: out = 12'h729;
            14'd 7234: out = 12'h72A;
            14'd 7235: out = 12'h72A;
            14'd 7236: out = 12'h72A;
            14'd 7237: out = 12'h72A;
            14'd 7238: out = 12'h72A;
            14'd 7239: out = 12'h72B;
            14'd 7240: out = 12'h72B;
            14'd 7241: out = 12'h72B;
            14'd 7242: out = 12'h72B;
            14'd 7243: out = 12'h72B;
            14'd 7244: out = 12'h72C;
            14'd 7245: out = 12'h72C;
            14'd 7246: out = 12'h72C;
            14'd 7247: out = 12'h72C;
            14'd 7248: out = 12'h72C;
            14'd 7249: out = 12'h72D;
            14'd 7250: out = 12'h72D;
            14'd 7251: out = 12'h72D;
            14'd 7252: out = 12'h72D;
            14'd 7253: out = 12'h72D;
            14'd 7254: out = 12'h72E;
            14'd 7255: out = 12'h72E;
            14'd 7256: out = 12'h72E;
            14'd 7257: out = 12'h72E;
            14'd 7258: out = 12'h72E;
            14'd 7259: out = 12'h72F;
            14'd 7260: out = 12'h72F;
            14'd 7261: out = 12'h72F;
            14'd 7262: out = 12'h72F;
            14'd 7263: out = 12'h72F;
            14'd 7264: out = 12'h730;
            14'd 7265: out = 12'h730;
            14'd 7266: out = 12'h730;
            14'd 7267: out = 12'h730;
            14'd 7268: out = 12'h730;
            14'd 7269: out = 12'h731;
            14'd 7270: out = 12'h731;
            14'd 7271: out = 12'h731;
            14'd 7272: out = 12'h731;
            14'd 7273: out = 12'h731;
            14'd 7274: out = 12'h732;
            14'd 7275: out = 12'h732;
            14'd 7276: out = 12'h732;
            14'd 7277: out = 12'h732;
            14'd 7278: out = 12'h732;
            14'd 7279: out = 12'h733;
            14'd 7280: out = 12'h733;
            14'd 7281: out = 12'h733;
            14'd 7282: out = 12'h733;
            14'd 7283: out = 12'h733;
            14'd 7284: out = 12'h734;
            14'd 7285: out = 12'h734;
            14'd 7286: out = 12'h734;
            14'd 7287: out = 12'h734;
            14'd 7288: out = 12'h734;
            14'd 7289: out = 12'h735;
            14'd 7290: out = 12'h735;
            14'd 7291: out = 12'h735;
            14'd 7292: out = 12'h735;
            14'd 7293: out = 12'h735;
            14'd 7294: out = 12'h736;
            14'd 7295: out = 12'h736;
            14'd 7296: out = 12'h736;
            14'd 7297: out = 12'h736;
            14'd 7298: out = 12'h736;
            14'd 7299: out = 12'h737;
            14'd 7300: out = 12'h737;
            14'd 7301: out = 12'h737;
            14'd 7302: out = 12'h737;
            14'd 7303: out = 12'h738;
            14'd 7304: out = 12'h738;
            14'd 7305: out = 12'h738;
            14'd 7306: out = 12'h738;
            14'd 7307: out = 12'h738;
            14'd 7308: out = 12'h739;
            14'd 7309: out = 12'h739;
            14'd 7310: out = 12'h739;
            14'd 7311: out = 12'h739;
            14'd 7312: out = 12'h739;
            14'd 7313: out = 12'h73A;
            14'd 7314: out = 12'h73A;
            14'd 7315: out = 12'h73A;
            14'd 7316: out = 12'h73A;
            14'd 7317: out = 12'h73A;
            14'd 7318: out = 12'h73B;
            14'd 7319: out = 12'h73B;
            14'd 7320: out = 12'h73B;
            14'd 7321: out = 12'h73B;
            14'd 7322: out = 12'h73B;
            14'd 7323: out = 12'h73C;
            14'd 7324: out = 12'h73C;
            14'd 7325: out = 12'h73C;
            14'd 7326: out = 12'h73C;
            14'd 7327: out = 12'h73C;
            14'd 7328: out = 12'h73D;
            14'd 7329: out = 12'h73D;
            14'd 7330: out = 12'h73D;
            14'd 7331: out = 12'h73D;
            14'd 7332: out = 12'h73D;
            14'd 7333: out = 12'h73E;
            14'd 7334: out = 12'h73E;
            14'd 7335: out = 12'h73E;
            14'd 7336: out = 12'h73E;
            14'd 7337: out = 12'h73E;
            14'd 7338: out = 12'h73F;
            14'd 7339: out = 12'h73F;
            14'd 7340: out = 12'h73F;
            14'd 7341: out = 12'h73F;
            14'd 7342: out = 12'h73F;
            14'd 7343: out = 12'h740;
            14'd 7344: out = 12'h740;
            14'd 7345: out = 12'h740;
            14'd 7346: out = 12'h740;
            14'd 7347: out = 12'h741;
            14'd 7348: out = 12'h741;
            14'd 7349: out = 12'h741;
            14'd 7350: out = 12'h741;
            14'd 7351: out = 12'h741;
            14'd 7352: out = 12'h742;
            14'd 7353: out = 12'h742;
            14'd 7354: out = 12'h742;
            14'd 7355: out = 12'h742;
            14'd 7356: out = 12'h742;
            14'd 7357: out = 12'h743;
            14'd 7358: out = 12'h743;
            14'd 7359: out = 12'h743;
            14'd 7360: out = 12'h743;
            14'd 7361: out = 12'h743;
            14'd 7362: out = 12'h744;
            14'd 7363: out = 12'h744;
            14'd 7364: out = 12'h744;
            14'd 7365: out = 12'h744;
            14'd 7366: out = 12'h744;
            14'd 7367: out = 12'h745;
            14'd 7368: out = 12'h745;
            14'd 7369: out = 12'h745;
            14'd 7370: out = 12'h745;
            14'd 7371: out = 12'h745;
            14'd 7372: out = 12'h746;
            14'd 7373: out = 12'h746;
            14'd 7374: out = 12'h746;
            14'd 7375: out = 12'h746;
            14'd 7376: out = 12'h746;
            14'd 7377: out = 12'h747;
            14'd 7378: out = 12'h747;
            14'd 7379: out = 12'h747;
            14'd 7380: out = 12'h747;
            14'd 7381: out = 12'h748;
            14'd 7382: out = 12'h748;
            14'd 7383: out = 12'h748;
            14'd 7384: out = 12'h748;
            14'd 7385: out = 12'h748;
            14'd 7386: out = 12'h749;
            14'd 7387: out = 12'h749;
            14'd 7388: out = 12'h749;
            14'd 7389: out = 12'h749;
            14'd 7390: out = 12'h749;
            14'd 7391: out = 12'h74A;
            14'd 7392: out = 12'h74A;
            14'd 7393: out = 12'h74A;
            14'd 7394: out = 12'h74A;
            14'd 7395: out = 12'h74A;
            14'd 7396: out = 12'h74B;
            14'd 7397: out = 12'h74B;
            14'd 7398: out = 12'h74B;
            14'd 7399: out = 12'h74B;
            14'd 7400: out = 12'h74B;
            14'd 7401: out = 12'h74C;
            14'd 7402: out = 12'h74C;
            14'd 7403: out = 12'h74C;
            14'd 7404: out = 12'h74C;
            14'd 7405: out = 12'h74C;
            14'd 7406: out = 12'h74D;
            14'd 7407: out = 12'h74D;
            14'd 7408: out = 12'h74D;
            14'd 7409: out = 12'h74D;
            14'd 7410: out = 12'h74E;
            14'd 7411: out = 12'h74E;
            14'd 7412: out = 12'h74E;
            14'd 7413: out = 12'h74E;
            14'd 7414: out = 12'h74E;
            14'd 7415: out = 12'h74F;
            14'd 7416: out = 12'h74F;
            14'd 7417: out = 12'h74F;
            14'd 7418: out = 12'h74F;
            14'd 7419: out = 12'h74F;
            14'd 7420: out = 12'h750;
            14'd 7421: out = 12'h750;
            14'd 7422: out = 12'h750;
            14'd 7423: out = 12'h750;
            14'd 7424: out = 12'h750;
            14'd 7425: out = 12'h751;
            14'd 7426: out = 12'h751;
            14'd 7427: out = 12'h751;
            14'd 7428: out = 12'h751;
            14'd 7429: out = 12'h752;
            14'd 7430: out = 12'h752;
            14'd 7431: out = 12'h752;
            14'd 7432: out = 12'h752;
            14'd 7433: out = 12'h752;
            14'd 7434: out = 12'h753;
            14'd 7435: out = 12'h753;
            14'd 7436: out = 12'h753;
            14'd 7437: out = 12'h753;
            14'd 7438: out = 12'h753;
            14'd 7439: out = 12'h754;
            14'd 7440: out = 12'h754;
            14'd 7441: out = 12'h754;
            14'd 7442: out = 12'h754;
            14'd 7443: out = 12'h754;
            14'd 7444: out = 12'h755;
            14'd 7445: out = 12'h755;
            14'd 7446: out = 12'h755;
            14'd 7447: out = 12'h755;
            14'd 7448: out = 12'h755;
            14'd 7449: out = 12'h756;
            14'd 7450: out = 12'h756;
            14'd 7451: out = 12'h756;
            14'd 7452: out = 12'h756;
            14'd 7453: out = 12'h757;
            14'd 7454: out = 12'h757;
            14'd 7455: out = 12'h757;
            14'd 7456: out = 12'h757;
            14'd 7457: out = 12'h757;
            14'd 7458: out = 12'h758;
            14'd 7459: out = 12'h758;
            14'd 7460: out = 12'h758;
            14'd 7461: out = 12'h758;
            14'd 7462: out = 12'h758;
            14'd 7463: out = 12'h759;
            14'd 7464: out = 12'h759;
            14'd 7465: out = 12'h759;
            14'd 7466: out = 12'h759;
            14'd 7467: out = 12'h759;
            14'd 7468: out = 12'h75A;
            14'd 7469: out = 12'h75A;
            14'd 7470: out = 12'h75A;
            14'd 7471: out = 12'h75A;
            14'd 7472: out = 12'h75B;
            14'd 7473: out = 12'h75B;
            14'd 7474: out = 12'h75B;
            14'd 7475: out = 12'h75B;
            14'd 7476: out = 12'h75B;
            14'd 7477: out = 12'h75C;
            14'd 7478: out = 12'h75C;
            14'd 7479: out = 12'h75C;
            14'd 7480: out = 12'h75C;
            14'd 7481: out = 12'h75C;
            14'd 7482: out = 12'h75D;
            14'd 7483: out = 12'h75D;
            14'd 7484: out = 12'h75D;
            14'd 7485: out = 12'h75D;
            14'd 7486: out = 12'h75E;
            14'd 7487: out = 12'h75E;
            14'd 7488: out = 12'h75E;
            14'd 7489: out = 12'h75E;
            14'd 7490: out = 12'h75E;
            14'd 7491: out = 12'h75F;
            14'd 7492: out = 12'h75F;
            14'd 7493: out = 12'h75F;
            14'd 7494: out = 12'h75F;
            14'd 7495: out = 12'h75F;
            14'd 7496: out = 12'h760;
            14'd 7497: out = 12'h760;
            14'd 7498: out = 12'h760;
            14'd 7499: out = 12'h760;
            14'd 7500: out = 12'h760;
            14'd 7501: out = 12'h761;
            14'd 7502: out = 12'h761;
            14'd 7503: out = 12'h761;
            14'd 7504: out = 12'h761;
            14'd 7505: out = 12'h762;
            14'd 7506: out = 12'h762;
            14'd 7507: out = 12'h762;
            14'd 7508: out = 12'h762;
            14'd 7509: out = 12'h762;
            14'd 7510: out = 12'h763;
            14'd 7511: out = 12'h763;
            14'd 7512: out = 12'h763;
            14'd 7513: out = 12'h763;
            14'd 7514: out = 12'h763;
            14'd 7515: out = 12'h764;
            14'd 7516: out = 12'h764;
            14'd 7517: out = 12'h764;
            14'd 7518: out = 12'h764;
            14'd 7519: out = 12'h765;
            14'd 7520: out = 12'h765;
            14'd 7521: out = 12'h765;
            14'd 7522: out = 12'h765;
            14'd 7523: out = 12'h765;
            14'd 7524: out = 12'h766;
            14'd 7525: out = 12'h766;
            14'd 7526: out = 12'h766;
            14'd 7527: out = 12'h766;
            14'd 7528: out = 12'h766;
            14'd 7529: out = 12'h767;
            14'd 7530: out = 12'h767;
            14'd 7531: out = 12'h767;
            14'd 7532: out = 12'h767;
            14'd 7533: out = 12'h768;
            14'd 7534: out = 12'h768;
            14'd 7535: out = 12'h768;
            14'd 7536: out = 12'h768;
            14'd 7537: out = 12'h768;
            14'd 7538: out = 12'h769;
            14'd 7539: out = 12'h769;
            14'd 7540: out = 12'h769;
            14'd 7541: out = 12'h769;
            14'd 7542: out = 12'h769;
            14'd 7543: out = 12'h76A;
            14'd 7544: out = 12'h76A;
            14'd 7545: out = 12'h76A;
            14'd 7546: out = 12'h76A;
            14'd 7547: out = 12'h76B;
            14'd 7548: out = 12'h76B;
            14'd 7549: out = 12'h76B;
            14'd 7550: out = 12'h76B;
            14'd 7551: out = 12'h76B;
            14'd 7552: out = 12'h76C;
            14'd 7553: out = 12'h76C;
            14'd 7554: out = 12'h76C;
            14'd 7555: out = 12'h76C;
            14'd 7556: out = 12'h76C;
            14'd 7557: out = 12'h76D;
            14'd 7558: out = 12'h76D;
            14'd 7559: out = 12'h76D;
            14'd 7560: out = 12'h76D;
            14'd 7561: out = 12'h76E;
            14'd 7562: out = 12'h76E;
            14'd 7563: out = 12'h76E;
            14'd 7564: out = 12'h76E;
            14'd 7565: out = 12'h76E;
            14'd 7566: out = 12'h76F;
            14'd 7567: out = 12'h76F;
            14'd 7568: out = 12'h76F;
            14'd 7569: out = 12'h76F;
            14'd 7570: out = 12'h76F;
            14'd 7571: out = 12'h770;
            14'd 7572: out = 12'h770;
            14'd 7573: out = 12'h770;
            14'd 7574: out = 12'h770;
            14'd 7575: out = 12'h771;
            14'd 7576: out = 12'h771;
            14'd 7577: out = 12'h771;
            14'd 7578: out = 12'h771;
            14'd 7579: out = 12'h771;
            14'd 7580: out = 12'h772;
            14'd 7581: out = 12'h772;
            14'd 7582: out = 12'h772;
            14'd 7583: out = 12'h772;
            14'd 7584: out = 12'h773;
            14'd 7585: out = 12'h773;
            14'd 7586: out = 12'h773;
            14'd 7587: out = 12'h773;
            14'd 7588: out = 12'h773;
            14'd 7589: out = 12'h774;
            14'd 7590: out = 12'h774;
            14'd 7591: out = 12'h774;
            14'd 7592: out = 12'h774;
            14'd 7593: out = 12'h774;
            14'd 7594: out = 12'h775;
            14'd 7595: out = 12'h775;
            14'd 7596: out = 12'h775;
            14'd 7597: out = 12'h775;
            14'd 7598: out = 12'h776;
            14'd 7599: out = 12'h776;
            14'd 7600: out = 12'h776;
            14'd 7601: out = 12'h776;
            14'd 7602: out = 12'h776;
            14'd 7603: out = 12'h777;
            14'd 7604: out = 12'h777;
            14'd 7605: out = 12'h777;
            14'd 7606: out = 12'h777;
            14'd 7607: out = 12'h777;
            14'd 7608: out = 12'h778;
            14'd 7609: out = 12'h778;
            14'd 7610: out = 12'h778;
            14'd 7611: out = 12'h778;
            14'd 7612: out = 12'h779;
            14'd 7613: out = 12'h779;
            14'd 7614: out = 12'h779;
            14'd 7615: out = 12'h779;
            14'd 7616: out = 12'h779;
            14'd 7617: out = 12'h77A;
            14'd 7618: out = 12'h77A;
            14'd 7619: out = 12'h77A;
            14'd 7620: out = 12'h77A;
            14'd 7621: out = 12'h77B;
            14'd 7622: out = 12'h77B;
            14'd 7623: out = 12'h77B;
            14'd 7624: out = 12'h77B;
            14'd 7625: out = 12'h77B;
            14'd 7626: out = 12'h77C;
            14'd 7627: out = 12'h77C;
            14'd 7628: out = 12'h77C;
            14'd 7629: out = 12'h77C;
            14'd 7630: out = 12'h77D;
            14'd 7631: out = 12'h77D;
            14'd 7632: out = 12'h77D;
            14'd 7633: out = 12'h77D;
            14'd 7634: out = 12'h77D;
            14'd 7635: out = 12'h77E;
            14'd 7636: out = 12'h77E;
            14'd 7637: out = 12'h77E;
            14'd 7638: out = 12'h77E;
            14'd 7639: out = 12'h77E;
            14'd 7640: out = 12'h77F;
            14'd 7641: out = 12'h77F;
            14'd 7642: out = 12'h77F;
            14'd 7643: out = 12'h77F;
            14'd 7644: out = 12'h780;
            14'd 7645: out = 12'h780;
            14'd 7646: out = 12'h780;
            14'd 7647: out = 12'h780;
            14'd 7648: out = 12'h780;
            14'd 7649: out = 12'h781;
            14'd 7650: out = 12'h781;
            14'd 7651: out = 12'h781;
            14'd 7652: out = 12'h781;
            14'd 7653: out = 12'h782;
            14'd 7654: out = 12'h782;
            14'd 7655: out = 12'h782;
            14'd 7656: out = 12'h782;
            14'd 7657: out = 12'h782;
            14'd 7658: out = 12'h783;
            14'd 7659: out = 12'h783;
            14'd 7660: out = 12'h783;
            14'd 7661: out = 12'h783;
            14'd 7662: out = 12'h784;
            14'd 7663: out = 12'h784;
            14'd 7664: out = 12'h784;
            14'd 7665: out = 12'h784;
            14'd 7666: out = 12'h784;
            14'd 7667: out = 12'h785;
            14'd 7668: out = 12'h785;
            14'd 7669: out = 12'h785;
            14'd 7670: out = 12'h785;
            14'd 7671: out = 12'h786;
            14'd 7672: out = 12'h786;
            14'd 7673: out = 12'h786;
            14'd 7674: out = 12'h786;
            14'd 7675: out = 12'h786;
            14'd 7676: out = 12'h787;
            14'd 7677: out = 12'h787;
            14'd 7678: out = 12'h787;
            14'd 7679: out = 12'h787;
            14'd 7680: out = 12'h788;
            14'd 7681: out = 12'h788;
            14'd 7682: out = 12'h788;
            14'd 7683: out = 12'h788;
            14'd 7684: out = 12'h788;
            14'd 7685: out = 12'h789;
            14'd 7686: out = 12'h789;
            14'd 7687: out = 12'h789;
            14'd 7688: out = 12'h789;
            14'd 7689: out = 12'h78A;
            14'd 7690: out = 12'h78A;
            14'd 7691: out = 12'h78A;
            14'd 7692: out = 12'h78A;
            14'd 7693: out = 12'h78A;
            14'd 7694: out = 12'h78B;
            14'd 7695: out = 12'h78B;
            14'd 7696: out = 12'h78B;
            14'd 7697: out = 12'h78B;
            14'd 7698: out = 12'h78C;
            14'd 7699: out = 12'h78C;
            14'd 7700: out = 12'h78C;
            14'd 7701: out = 12'h78C;
            14'd 7702: out = 12'h78C;
            14'd 7703: out = 12'h78D;
            14'd 7704: out = 12'h78D;
            14'd 7705: out = 12'h78D;
            14'd 7706: out = 12'h78D;
            14'd 7707: out = 12'h78E;
            14'd 7708: out = 12'h78E;
            14'd 7709: out = 12'h78E;
            14'd 7710: out = 12'h78E;
            14'd 7711: out = 12'h78E;
            14'd 7712: out = 12'h78F;
            14'd 7713: out = 12'h78F;
            14'd 7714: out = 12'h78F;
            14'd 7715: out = 12'h78F;
            14'd 7716: out = 12'h790;
            14'd 7717: out = 12'h790;
            14'd 7718: out = 12'h790;
            14'd 7719: out = 12'h790;
            14'd 7720: out = 12'h790;
            14'd 7721: out = 12'h791;
            14'd 7722: out = 12'h791;
            14'd 7723: out = 12'h791;
            14'd 7724: out = 12'h791;
            14'd 7725: out = 12'h792;
            14'd 7726: out = 12'h792;
            14'd 7727: out = 12'h792;
            14'd 7728: out = 12'h792;
            14'd 7729: out = 12'h792;
            14'd 7730: out = 12'h793;
            14'd 7731: out = 12'h793;
            14'd 7732: out = 12'h793;
            14'd 7733: out = 12'h793;
            14'd 7734: out = 12'h794;
            14'd 7735: out = 12'h794;
            14'd 7736: out = 12'h794;
            14'd 7737: out = 12'h794;
            14'd 7738: out = 12'h794;
            14'd 7739: out = 12'h795;
            14'd 7740: out = 12'h795;
            14'd 7741: out = 12'h795;
            14'd 7742: out = 12'h795;
            14'd 7743: out = 12'h796;
            14'd 7744: out = 12'h796;
            14'd 7745: out = 12'h796;
            14'd 7746: out = 12'h796;
            14'd 7747: out = 12'h796;
            14'd 7748: out = 12'h797;
            14'd 7749: out = 12'h797;
            14'd 7750: out = 12'h797;
            14'd 7751: out = 12'h797;
            14'd 7752: out = 12'h798;
            14'd 7753: out = 12'h798;
            14'd 7754: out = 12'h798;
            14'd 7755: out = 12'h798;
            14'd 7756: out = 12'h799;
            14'd 7757: out = 12'h799;
            14'd 7758: out = 12'h799;
            14'd 7759: out = 12'h799;
            14'd 7760: out = 12'h799;
            14'd 7761: out = 12'h79A;
            14'd 7762: out = 12'h79A;
            14'd 7763: out = 12'h79A;
            14'd 7764: out = 12'h79A;
            14'd 7765: out = 12'h79B;
            14'd 7766: out = 12'h79B;
            14'd 7767: out = 12'h79B;
            14'd 7768: out = 12'h79B;
            14'd 7769: out = 12'h79B;
            14'd 7770: out = 12'h79C;
            14'd 7771: out = 12'h79C;
            14'd 7772: out = 12'h79C;
            14'd 7773: out = 12'h79C;
            14'd 7774: out = 12'h79D;
            14'd 7775: out = 12'h79D;
            14'd 7776: out = 12'h79D;
            14'd 7777: out = 12'h79D;
            14'd 7778: out = 12'h79D;
            14'd 7779: out = 12'h79E;
            14'd 7780: out = 12'h79E;
            14'd 7781: out = 12'h79E;
            14'd 7782: out = 12'h79E;
            14'd 7783: out = 12'h79F;
            14'd 7784: out = 12'h79F;
            14'd 7785: out = 12'h79F;
            14'd 7786: out = 12'h79F;
            14'd 7787: out = 12'h7A0;
            14'd 7788: out = 12'h7A0;
            14'd 7789: out = 12'h7A0;
            14'd 7790: out = 12'h7A0;
            14'd 7791: out = 12'h7A0;
            14'd 7792: out = 12'h7A1;
            14'd 7793: out = 12'h7A1;
            14'd 7794: out = 12'h7A1;
            14'd 7795: out = 12'h7A1;
            14'd 7796: out = 12'h7A2;
            14'd 7797: out = 12'h7A2;
            14'd 7798: out = 12'h7A2;
            14'd 7799: out = 12'h7A2;
            14'd 7800: out = 12'h7A2;
            14'd 7801: out = 12'h7A3;
            14'd 7802: out = 12'h7A3;
            14'd 7803: out = 12'h7A3;
            14'd 7804: out = 12'h7A3;
            14'd 7805: out = 12'h7A4;
            14'd 7806: out = 12'h7A4;
            14'd 7807: out = 12'h7A4;
            14'd 7808: out = 12'h7A4;
            14'd 7809: out = 12'h7A5;
            14'd 7810: out = 12'h7A5;
            14'd 7811: out = 12'h7A5;
            14'd 7812: out = 12'h7A5;
            14'd 7813: out = 12'h7A5;
            14'd 7814: out = 12'h7A6;
            14'd 7815: out = 12'h7A6;
            14'd 7816: out = 12'h7A6;
            14'd 7817: out = 12'h7A6;
            14'd 7818: out = 12'h7A7;
            14'd 7819: out = 12'h7A7;
            14'd 7820: out = 12'h7A7;
            14'd 7821: out = 12'h7A7;
            14'd 7822: out = 12'h7A7;
            14'd 7823: out = 12'h7A8;
            14'd 7824: out = 12'h7A8;
            14'd 7825: out = 12'h7A8;
            14'd 7826: out = 12'h7A8;
            14'd 7827: out = 12'h7A9;
            14'd 7828: out = 12'h7A9;
            14'd 7829: out = 12'h7A9;
            14'd 7830: out = 12'h7A9;
            14'd 7831: out = 12'h7AA;
            14'd 7832: out = 12'h7AA;
            14'd 7833: out = 12'h7AA;
            14'd 7834: out = 12'h7AA;
            14'd 7835: out = 12'h7AA;
            14'd 7836: out = 12'h7AB;
            14'd 7837: out = 12'h7AB;
            14'd 7838: out = 12'h7AB;
            14'd 7839: out = 12'h7AB;
            14'd 7840: out = 12'h7AC;
            14'd 7841: out = 12'h7AC;
            14'd 7842: out = 12'h7AC;
            14'd 7843: out = 12'h7AC;
            14'd 7844: out = 12'h7AD;
            14'd 7845: out = 12'h7AD;
            14'd 7846: out = 12'h7AD;
            14'd 7847: out = 12'h7AD;
            14'd 7848: out = 12'h7AD;
            14'd 7849: out = 12'h7AE;
            14'd 7850: out = 12'h7AE;
            14'd 7851: out = 12'h7AE;
            14'd 7852: out = 12'h7AE;
            14'd 7853: out = 12'h7AF;
            14'd 7854: out = 12'h7AF;
            14'd 7855: out = 12'h7AF;
            14'd 7856: out = 12'h7AF;
            14'd 7857: out = 12'h7B0;
            14'd 7858: out = 12'h7B0;
            14'd 7859: out = 12'h7B0;
            14'd 7860: out = 12'h7B0;
            14'd 7861: out = 12'h7B0;
            14'd 7862: out = 12'h7B1;
            14'd 7863: out = 12'h7B1;
            14'd 7864: out = 12'h7B1;
            14'd 7865: out = 12'h7B1;
            14'd 7866: out = 12'h7B2;
            14'd 7867: out = 12'h7B2;
            14'd 7868: out = 12'h7B2;
            14'd 7869: out = 12'h7B2;
            14'd 7870: out = 12'h7B3;
            14'd 7871: out = 12'h7B3;
            14'd 7872: out = 12'h7B3;
            14'd 7873: out = 12'h7B3;
            14'd 7874: out = 12'h7B3;
            14'd 7875: out = 12'h7B4;
            14'd 7876: out = 12'h7B4;
            14'd 7877: out = 12'h7B4;
            14'd 7878: out = 12'h7B4;
            14'd 7879: out = 12'h7B5;
            14'd 7880: out = 12'h7B5;
            14'd 7881: out = 12'h7B5;
            14'd 7882: out = 12'h7B5;
            14'd 7883: out = 12'h7B6;
            14'd 7884: out = 12'h7B6;
            14'd 7885: out = 12'h7B6;
            14'd 7886: out = 12'h7B6;
            14'd 7887: out = 12'h7B6;
            14'd 7888: out = 12'h7B7;
            14'd 7889: out = 12'h7B7;
            14'd 7890: out = 12'h7B7;
            14'd 7891: out = 12'h7B7;
            14'd 7892: out = 12'h7B8;
            14'd 7893: out = 12'h7B8;
            14'd 7894: out = 12'h7B8;
            14'd 7895: out = 12'h7B8;
            14'd 7896: out = 12'h7B9;
            14'd 7897: out = 12'h7B9;
            14'd 7898: out = 12'h7B9;
            14'd 7899: out = 12'h7B9;
            14'd 7900: out = 12'h7BA;
            14'd 7901: out = 12'h7BA;
            14'd 7902: out = 12'h7BA;
            14'd 7903: out = 12'h7BA;
            14'd 7904: out = 12'h7BA;
            14'd 7905: out = 12'h7BB;
            14'd 7906: out = 12'h7BB;
            14'd 7907: out = 12'h7BB;
            14'd 7908: out = 12'h7BB;
            14'd 7909: out = 12'h7BC;
            14'd 7910: out = 12'h7BC;
            14'd 7911: out = 12'h7BC;
            14'd 7912: out = 12'h7BC;
            14'd 7913: out = 12'h7BD;
            14'd 7914: out = 12'h7BD;
            14'd 7915: out = 12'h7BD;
            14'd 7916: out = 12'h7BD;
            14'd 7917: out = 12'h7BD;
            14'd 7918: out = 12'h7BE;
            14'd 7919: out = 12'h7BE;
            14'd 7920: out = 12'h7BE;
            14'd 7921: out = 12'h7BE;
            14'd 7922: out = 12'h7BF;
            14'd 7923: out = 12'h7BF;
            14'd 7924: out = 12'h7BF;
            14'd 7925: out = 12'h7BF;
            14'd 7926: out = 12'h7C0;
            14'd 7927: out = 12'h7C0;
            14'd 7928: out = 12'h7C0;
            14'd 7929: out = 12'h7C0;
            14'd 7930: out = 12'h7C1;
            14'd 7931: out = 12'h7C1;
            14'd 7932: out = 12'h7C1;
            14'd 7933: out = 12'h7C1;
            14'd 7934: out = 12'h7C1;
            14'd 7935: out = 12'h7C2;
            14'd 7936: out = 12'h7C2;
            14'd 7937: out = 12'h7C2;
            14'd 7938: out = 12'h7C2;
            14'd 7939: out = 12'h7C3;
            14'd 7940: out = 12'h7C3;
            14'd 7941: out = 12'h7C3;
            14'd 7942: out = 12'h7C3;
            14'd 7943: out = 12'h7C4;
            14'd 7944: out = 12'h7C4;
            14'd 7945: out = 12'h7C4;
            14'd 7946: out = 12'h7C4;
            14'd 7947: out = 12'h7C5;
            14'd 7948: out = 12'h7C5;
            14'd 7949: out = 12'h7C5;
            14'd 7950: out = 12'h7C5;
            14'd 7951: out = 12'h7C5;
            14'd 7952: out = 12'h7C6;
            14'd 7953: out = 12'h7C6;
            14'd 7954: out = 12'h7C6;
            14'd 7955: out = 12'h7C6;
            14'd 7956: out = 12'h7C7;
            14'd 7957: out = 12'h7C7;
            14'd 7958: out = 12'h7C7;
            14'd 7959: out = 12'h7C7;
            14'd 7960: out = 12'h7C8;
            14'd 7961: out = 12'h7C8;
            14'd 7962: out = 12'h7C8;
            14'd 7963: out = 12'h7C8;
            14'd 7964: out = 12'h7C9;
            14'd 7965: out = 12'h7C9;
            14'd 7966: out = 12'h7C9;
            14'd 7967: out = 12'h7C9;
            14'd 7968: out = 12'h7C9;
            14'd 7969: out = 12'h7CA;
            14'd 7970: out = 12'h7CA;
            14'd 7971: out = 12'h7CA;
            14'd 7972: out = 12'h7CA;
            14'd 7973: out = 12'h7CB;
            14'd 7974: out = 12'h7CB;
            14'd 7975: out = 12'h7CB;
            14'd 7976: out = 12'h7CB;
            14'd 7977: out = 12'h7CC;
            14'd 7978: out = 12'h7CC;
            14'd 7979: out = 12'h7CC;
            14'd 7980: out = 12'h7CC;
            14'd 7981: out = 12'h7CD;
            14'd 7982: out = 12'h7CD;
            14'd 7983: out = 12'h7CD;
            14'd 7984: out = 12'h7CD;
            14'd 7985: out = 12'h7CE;
            14'd 7986: out = 12'h7CE;
            14'd 7987: out = 12'h7CE;
            14'd 7988: out = 12'h7CE;
            14'd 7989: out = 12'h7CE;
            14'd 7990: out = 12'h7CF;
            14'd 7991: out = 12'h7CF;
            14'd 7992: out = 12'h7CF;
            14'd 7993: out = 12'h7CF;
            14'd 7994: out = 12'h7D0;
            14'd 7995: out = 12'h7D0;
            14'd 7996: out = 12'h7D0;
            14'd 7997: out = 12'h7D0;
            14'd 7998: out = 12'h7D1;
            14'd 7999: out = 12'h7D1;
            14'd 8000: out = 12'h7D1;
            14'd 8001: out = 12'h7D1;
            14'd 8002: out = 12'h7D2;
            14'd 8003: out = 12'h7D2;
            14'd 8004: out = 12'h7D2;
            14'd 8005: out = 12'h7D2;
            14'd 8006: out = 12'h7D3;
            14'd 8007: out = 12'h7D3;
            14'd 8008: out = 12'h7D3;
            14'd 8009: out = 12'h7D3;
            14'd 8010: out = 12'h7D3;
            14'd 8011: out = 12'h7D4;
            14'd 8012: out = 12'h7D4;
            14'd 8013: out = 12'h7D4;
            14'd 8014: out = 12'h7D4;
            14'd 8015: out = 12'h7D5;
            14'd 8016: out = 12'h7D5;
            14'd 8017: out = 12'h7D5;
            14'd 8018: out = 12'h7D5;
            14'd 8019: out = 12'h7D6;
            14'd 8020: out = 12'h7D6;
            14'd 8021: out = 12'h7D6;
            14'd 8022: out = 12'h7D6;
            14'd 8023: out = 12'h7D7;
            14'd 8024: out = 12'h7D7;
            14'd 8025: out = 12'h7D7;
            14'd 8026: out = 12'h7D7;
            14'd 8027: out = 12'h7D8;
            14'd 8028: out = 12'h7D8;
            14'd 8029: out = 12'h7D8;
            14'd 8030: out = 12'h7D8;
            14'd 8031: out = 12'h7D9;
            14'd 8032: out = 12'h7D9;
            14'd 8033: out = 12'h7D9;
            14'd 8034: out = 12'h7D9;
            14'd 8035: out = 12'h7D9;
            14'd 8036: out = 12'h7DA;
            14'd 8037: out = 12'h7DA;
            14'd 8038: out = 12'h7DA;
            14'd 8039: out = 12'h7DA;
            14'd 8040: out = 12'h7DB;
            14'd 8041: out = 12'h7DB;
            14'd 8042: out = 12'h7DB;
            14'd 8043: out = 12'h7DB;
            14'd 8044: out = 12'h7DC;
            14'd 8045: out = 12'h7DC;
            14'd 8046: out = 12'h7DC;
            14'd 8047: out = 12'h7DC;
            14'd 8048: out = 12'h7DD;
            14'd 8049: out = 12'h7DD;
            14'd 8050: out = 12'h7DD;
            14'd 8051: out = 12'h7DD;
            14'd 8052: out = 12'h7DE;
            14'd 8053: out = 12'h7DE;
            14'd 8054: out = 12'h7DE;
            14'd 8055: out = 12'h7DE;
            14'd 8056: out = 12'h7DF;
            14'd 8057: out = 12'h7DF;
            14'd 8058: out = 12'h7DF;
            14'd 8059: out = 12'h7DF;
            14'd 8060: out = 12'h7E0;
            14'd 8061: out = 12'h7E0;
            14'd 8062: out = 12'h7E0;
            14'd 8063: out = 12'h7E0;
            14'd 8064: out = 12'h7E0;
            14'd 8065: out = 12'h7E1;
            14'd 8066: out = 12'h7E1;
            14'd 8067: out = 12'h7E1;
            14'd 8068: out = 12'h7E1;
            14'd 8069: out = 12'h7E2;
            14'd 8070: out = 12'h7E2;
            14'd 8071: out = 12'h7E2;
            14'd 8072: out = 12'h7E2;
            14'd 8073: out = 12'h7E3;
            14'd 8074: out = 12'h7E3;
            14'd 8075: out = 12'h7E3;
            14'd 8076: out = 12'h7E3;
            14'd 8077: out = 12'h7E4;
            14'd 8078: out = 12'h7E4;
            14'd 8079: out = 12'h7E4;
            14'd 8080: out = 12'h7E4;
            14'd 8081: out = 12'h7E5;
            14'd 8082: out = 12'h7E5;
            14'd 8083: out = 12'h7E5;
            14'd 8084: out = 12'h7E5;
            14'd 8085: out = 12'h7E6;
            14'd 8086: out = 12'h7E6;
            14'd 8087: out = 12'h7E6;
            14'd 8088: out = 12'h7E6;
            14'd 8089: out = 12'h7E7;
            14'd 8090: out = 12'h7E7;
            14'd 8091: out = 12'h7E7;
            14'd 8092: out = 12'h7E7;
            14'd 8093: out = 12'h7E8;
            14'd 8094: out = 12'h7E8;
            14'd 8095: out = 12'h7E8;
            14'd 8096: out = 12'h7E8;
            14'd 8097: out = 12'h7E9;
            14'd 8098: out = 12'h7E9;
            14'd 8099: out = 12'h7E9;
            14'd 8100: out = 12'h7E9;
            14'd 8101: out = 12'h7E9;
            14'd 8102: out = 12'h7EA;
            14'd 8103: out = 12'h7EA;
            14'd 8104: out = 12'h7EA;
            14'd 8105: out = 12'h7EA;
            14'd 8106: out = 12'h7EB;
            14'd 8107: out = 12'h7EB;
            14'd 8108: out = 12'h7EB;
            14'd 8109: out = 12'h7EB;
            14'd 8110: out = 12'h7EC;
            14'd 8111: out = 12'h7EC;
            14'd 8112: out = 12'h7EC;
            14'd 8113: out = 12'h7EC;
            14'd 8114: out = 12'h7ED;
            14'd 8115: out = 12'h7ED;
            14'd 8116: out = 12'h7ED;
            14'd 8117: out = 12'h7ED;
            14'd 8118: out = 12'h7EE;
            14'd 8119: out = 12'h7EE;
            14'd 8120: out = 12'h7EE;
            14'd 8121: out = 12'h7EE;
            14'd 8122: out = 12'h7EF;
            14'd 8123: out = 12'h7EF;
            14'd 8124: out = 12'h7EF;
            14'd 8125: out = 12'h7EF;
            14'd 8126: out = 12'h7F0;
            14'd 8127: out = 12'h7F0;
            14'd 8128: out = 12'h7F0;
            14'd 8129: out = 12'h7F0;
            14'd 8130: out = 12'h7F1;
            14'd 8131: out = 12'h7F1;
            14'd 8132: out = 12'h7F1;
            14'd 8133: out = 12'h7F1;
            14'd 8134: out = 12'h7F2;
            14'd 8135: out = 12'h7F2;
            14'd 8136: out = 12'h7F2;
            14'd 8137: out = 12'h7F2;
            14'd 8138: out = 12'h7F3;
            14'd 8139: out = 12'h7F3;
            14'd 8140: out = 12'h7F3;
            14'd 8141: out = 12'h7F3;
            14'd 8142: out = 12'h7F4;
            14'd 8143: out = 12'h7F4;
            14'd 8144: out = 12'h7F4;
            14'd 8145: out = 12'h7F4;
            14'd 8146: out = 12'h7F5;
            14'd 8147: out = 12'h7F5;
            14'd 8148: out = 12'h7F5;
            14'd 8149: out = 12'h7F5;
            14'd 8150: out = 12'h7F6;
            14'd 8151: out = 12'h7F6;
            14'd 8152: out = 12'h7F6;
            14'd 8153: out = 12'h7F6;
            14'd 8154: out = 12'h7F7;
            14'd 8155: out = 12'h7F7;
            14'd 8156: out = 12'h7F7;
            14'd 8157: out = 12'h7F7;
            14'd 8158: out = 12'h7F8;
            14'd 8159: out = 12'h7F8;
            14'd 8160: out = 12'h7F8;
            14'd 8161: out = 12'h7F8;
            14'd 8162: out = 12'h7F9;
            14'd 8163: out = 12'h7F9;
            14'd 8164: out = 12'h7F9;
            14'd 8165: out = 12'h7F9;
            14'd 8166: out = 12'h7FA;
            14'd 8167: out = 12'h7FA;
            14'd 8168: out = 12'h7FA;
            14'd 8169: out = 12'h7FA;
            14'd 8170: out = 12'h7FB;
            14'd 8171: out = 12'h7FB;
            14'd 8172: out = 12'h7FB;
            14'd 8173: out = 12'h7FB;
            14'd 8174: out = 12'h7FC;
            14'd 8175: out = 12'h7FC;
            14'd 8176: out = 12'h7FC;
            14'd 8177: out = 12'h7FC;
            14'd 8178: out = 12'h7FD;
            14'd 8179: out = 12'h7FD;
            14'd 8180: out = 12'h7FD;
            14'd 8181: out = 12'h7FD;
            14'd 8182: out = 12'h7FE;
            14'd 8183: out = 12'h7FE;
            14'd 8184: out = 12'h7FE;
            14'd 8185: out = 12'h7FE;
            14'd 8186: out = 12'h7FF;
            14'd 8187: out = 12'h7FF;
            14'd 8188: out = 12'h7FF;
            14'd 8189: out = 12'h7FF;
            14'd 8190: out = 12'h800;
            14'd 8191: out = 12'h800;
            14'd 8192: out = 12'h800;
            14'd 8193: out = 12'h800;
            14'd 8194: out = 12'h801;
            14'd 8195: out = 12'h801;
            14'd 8196: out = 12'h801;
            14'd 8197: out = 12'h801;
            14'd 8198: out = 12'h802;
            14'd 8199: out = 12'h802;
            14'd 8200: out = 12'h802;
            14'd 8201: out = 12'h802;
            14'd 8202: out = 12'h803;
            14'd 8203: out = 12'h803;
            14'd 8204: out = 12'h803;
            14'd 8205: out = 12'h803;
            14'd 8206: out = 12'h804;
            14'd 8207: out = 12'h804;
            14'd 8208: out = 12'h804;
            14'd 8209: out = 12'h804;
            14'd 8210: out = 12'h805;
            14'd 8211: out = 12'h805;
            14'd 8212: out = 12'h805;
            14'd 8213: out = 12'h805;
            14'd 8214: out = 12'h806;
            14'd 8215: out = 12'h806;
            14'd 8216: out = 12'h806;
            14'd 8217: out = 12'h806;
            14'd 8218: out = 12'h807;
            14'd 8219: out = 12'h807;
            14'd 8220: out = 12'h807;
            14'd 8221: out = 12'h807;
            14'd 8222: out = 12'h808;
            14'd 8223: out = 12'h808;
            14'd 8224: out = 12'h808;
            14'd 8225: out = 12'h808;
            14'd 8226: out = 12'h809;
            14'd 8227: out = 12'h809;
            14'd 8228: out = 12'h809;
            14'd 8229: out = 12'h809;
            14'd 8230: out = 12'h80A;
            14'd 8231: out = 12'h80A;
            14'd 8232: out = 12'h80A;
            14'd 8233: out = 12'h80A;
            14'd 8234: out = 12'h80B;
            14'd 8235: out = 12'h80B;
            14'd 8236: out = 12'h80B;
            14'd 8237: out = 12'h80B;
            14'd 8238: out = 12'h80C;
            14'd 8239: out = 12'h80C;
            14'd 8240: out = 12'h80C;
            14'd 8241: out = 12'h80C;
            14'd 8242: out = 12'h80D;
            14'd 8243: out = 12'h80D;
            14'd 8244: out = 12'h80D;
            14'd 8245: out = 12'h80D;
            14'd 8246: out = 12'h80E;
            14'd 8247: out = 12'h80E;
            14'd 8248: out = 12'h80E;
            14'd 8249: out = 12'h80E;
            14'd 8250: out = 12'h80F;
            14'd 8251: out = 12'h80F;
            14'd 8252: out = 12'h80F;
            14'd 8253: out = 12'h80F;
            14'd 8254: out = 12'h810;
            14'd 8255: out = 12'h810;
            14'd 8256: out = 12'h810;
            14'd 8257: out = 12'h810;
            14'd 8258: out = 12'h811;
            14'd 8259: out = 12'h811;
            14'd 8260: out = 12'h811;
            14'd 8261: out = 12'h811;
            14'd 8262: out = 12'h812;
            14'd 8263: out = 12'h812;
            14'd 8264: out = 12'h812;
            14'd 8265: out = 12'h812;
            14'd 8266: out = 12'h813;
            14'd 8267: out = 12'h813;
            14'd 8268: out = 12'h813;
            14'd 8269: out = 12'h813;
            14'd 8270: out = 12'h814;
            14'd 8271: out = 12'h814;
            14'd 8272: out = 12'h814;
            14'd 8273: out = 12'h814;
            14'd 8274: out = 12'h815;
            14'd 8275: out = 12'h815;
            14'd 8276: out = 12'h815;
            14'd 8277: out = 12'h815;
            14'd 8278: out = 12'h816;
            14'd 8279: out = 12'h816;
            14'd 8280: out = 12'h816;
            14'd 8281: out = 12'h816;
            14'd 8282: out = 12'h817;
            14'd 8283: out = 12'h817;
            14'd 8284: out = 12'h817;
            14'd 8285: out = 12'h818;
            14'd 8286: out = 12'h818;
            14'd 8287: out = 12'h818;
            14'd 8288: out = 12'h818;
            14'd 8289: out = 12'h819;
            14'd 8290: out = 12'h819;
            14'd 8291: out = 12'h819;
            14'd 8292: out = 12'h819;
            14'd 8293: out = 12'h81A;
            14'd 8294: out = 12'h81A;
            14'd 8295: out = 12'h81A;
            14'd 8296: out = 12'h81A;
            14'd 8297: out = 12'h81B;
            14'd 8298: out = 12'h81B;
            14'd 8299: out = 12'h81B;
            14'd 8300: out = 12'h81B;
            14'd 8301: out = 12'h81C;
            14'd 8302: out = 12'h81C;
            14'd 8303: out = 12'h81C;
            14'd 8304: out = 12'h81C;
            14'd 8305: out = 12'h81D;
            14'd 8306: out = 12'h81D;
            14'd 8307: out = 12'h81D;
            14'd 8308: out = 12'h81D;
            14'd 8309: out = 12'h81E;
            14'd 8310: out = 12'h81E;
            14'd 8311: out = 12'h81E;
            14'd 8312: out = 12'h81E;
            14'd 8313: out = 12'h81F;
            14'd 8314: out = 12'h81F;
            14'd 8315: out = 12'h81F;
            14'd 8316: out = 12'h81F;
            14'd 8317: out = 12'h820;
            14'd 8318: out = 12'h820;
            14'd 8319: out = 12'h820;
            14'd 8320: out = 12'h821;
            14'd 8321: out = 12'h821;
            14'd 8322: out = 12'h821;
            14'd 8323: out = 12'h821;
            14'd 8324: out = 12'h822;
            14'd 8325: out = 12'h822;
            14'd 8326: out = 12'h822;
            14'd 8327: out = 12'h822;
            14'd 8328: out = 12'h823;
            14'd 8329: out = 12'h823;
            14'd 8330: out = 12'h823;
            14'd 8331: out = 12'h823;
            14'd 8332: out = 12'h824;
            14'd 8333: out = 12'h824;
            14'd 8334: out = 12'h824;
            14'd 8335: out = 12'h824;
            14'd 8336: out = 12'h825;
            14'd 8337: out = 12'h825;
            14'd 8338: out = 12'h825;
            14'd 8339: out = 12'h825;
            14'd 8340: out = 12'h826;
            14'd 8341: out = 12'h826;
            14'd 8342: out = 12'h826;
            14'd 8343: out = 12'h826;
            14'd 8344: out = 12'h827;
            14'd 8345: out = 12'h827;
            14'd 8346: out = 12'h827;
            14'd 8347: out = 12'h827;
            14'd 8348: out = 12'h828;
            14'd 8349: out = 12'h828;
            14'd 8350: out = 12'h828;
            14'd 8351: out = 12'h829;
            14'd 8352: out = 12'h829;
            14'd 8353: out = 12'h829;
            14'd 8354: out = 12'h829;
            14'd 8355: out = 12'h82A;
            14'd 8356: out = 12'h82A;
            14'd 8357: out = 12'h82A;
            14'd 8358: out = 12'h82A;
            14'd 8359: out = 12'h82B;
            14'd 8360: out = 12'h82B;
            14'd 8361: out = 12'h82B;
            14'd 8362: out = 12'h82B;
            14'd 8363: out = 12'h82C;
            14'd 8364: out = 12'h82C;
            14'd 8365: out = 12'h82C;
            14'd 8366: out = 12'h82C;
            14'd 8367: out = 12'h82D;
            14'd 8368: out = 12'h82D;
            14'd 8369: out = 12'h82D;
            14'd 8370: out = 12'h82D;
            14'd 8371: out = 12'h82E;
            14'd 8372: out = 12'h82E;
            14'd 8373: out = 12'h82E;
            14'd 8374: out = 12'h82F;
            14'd 8375: out = 12'h82F;
            14'd 8376: out = 12'h82F;
            14'd 8377: out = 12'h82F;
            14'd 8378: out = 12'h830;
            14'd 8379: out = 12'h830;
            14'd 8380: out = 12'h830;
            14'd 8381: out = 12'h830;
            14'd 8382: out = 12'h831;
            14'd 8383: out = 12'h831;
            14'd 8384: out = 12'h831;
            14'd 8385: out = 12'h831;
            14'd 8386: out = 12'h832;
            14'd 8387: out = 12'h832;
            14'd 8388: out = 12'h832;
            14'd 8389: out = 12'h832;
            14'd 8390: out = 12'h833;
            14'd 8391: out = 12'h833;
            14'd 8392: out = 12'h833;
            14'd 8393: out = 12'h834;
            14'd 8394: out = 12'h834;
            14'd 8395: out = 12'h834;
            14'd 8396: out = 12'h834;
            14'd 8397: out = 12'h835;
            14'd 8398: out = 12'h835;
            14'd 8399: out = 12'h835;
            14'd 8400: out = 12'h835;
            14'd 8401: out = 12'h836;
            14'd 8402: out = 12'h836;
            14'd 8403: out = 12'h836;
            14'd 8404: out = 12'h836;
            14'd 8405: out = 12'h837;
            14'd 8406: out = 12'h837;
            14'd 8407: out = 12'h837;
            14'd 8408: out = 12'h837;
            14'd 8409: out = 12'h838;
            14'd 8410: out = 12'h838;
            14'd 8411: out = 12'h838;
            14'd 8412: out = 12'h839;
            14'd 8413: out = 12'h839;
            14'd 8414: out = 12'h839;
            14'd 8415: out = 12'h839;
            14'd 8416: out = 12'h83A;
            14'd 8417: out = 12'h83A;
            14'd 8418: out = 12'h83A;
            14'd 8419: out = 12'h83A;
            14'd 8420: out = 12'h83B;
            14'd 8421: out = 12'h83B;
            14'd 8422: out = 12'h83B;
            14'd 8423: out = 12'h83B;
            14'd 8424: out = 12'h83C;
            14'd 8425: out = 12'h83C;
            14'd 8426: out = 12'h83C;
            14'd 8427: out = 12'h83C;
            14'd 8428: out = 12'h83D;
            14'd 8429: out = 12'h83D;
            14'd 8430: out = 12'h83D;
            14'd 8431: out = 12'h83E;
            14'd 8432: out = 12'h83E;
            14'd 8433: out = 12'h83E;
            14'd 8434: out = 12'h83E;
            14'd 8435: out = 12'h83F;
            14'd 8436: out = 12'h83F;
            14'd 8437: out = 12'h83F;
            14'd 8438: out = 12'h83F;
            14'd 8439: out = 12'h840;
            14'd 8440: out = 12'h840;
            14'd 8441: out = 12'h840;
            14'd 8442: out = 12'h840;
            14'd 8443: out = 12'h841;
            14'd 8444: out = 12'h841;
            14'd 8445: out = 12'h841;
            14'd 8446: out = 12'h842;
            14'd 8447: out = 12'h842;
            14'd 8448: out = 12'h842;
            14'd 8449: out = 12'h842;
            14'd 8450: out = 12'h843;
            14'd 8451: out = 12'h843;
            14'd 8452: out = 12'h843;
            14'd 8453: out = 12'h843;
            14'd 8454: out = 12'h844;
            14'd 8455: out = 12'h844;
            14'd 8456: out = 12'h844;
            14'd 8457: out = 12'h844;
            14'd 8458: out = 12'h845;
            14'd 8459: out = 12'h845;
            14'd 8460: out = 12'h845;
            14'd 8461: out = 12'h846;
            14'd 8462: out = 12'h846;
            14'd 8463: out = 12'h846;
            14'd 8464: out = 12'h846;
            14'd 8465: out = 12'h847;
            14'd 8466: out = 12'h847;
            14'd 8467: out = 12'h847;
            14'd 8468: out = 12'h847;
            14'd 8469: out = 12'h848;
            14'd 8470: out = 12'h848;
            14'd 8471: out = 12'h848;
            14'd 8472: out = 12'h848;
            14'd 8473: out = 12'h849;
            14'd 8474: out = 12'h849;
            14'd 8475: out = 12'h849;
            14'd 8476: out = 12'h84A;
            14'd 8477: out = 12'h84A;
            14'd 8478: out = 12'h84A;
            14'd 8479: out = 12'h84A;
            14'd 8480: out = 12'h84B;
            14'd 8481: out = 12'h84B;
            14'd 8482: out = 12'h84B;
            14'd 8483: out = 12'h84B;
            14'd 8484: out = 12'h84C;
            14'd 8485: out = 12'h84C;
            14'd 8486: out = 12'h84C;
            14'd 8487: out = 12'h84D;
            14'd 8488: out = 12'h84D;
            14'd 8489: out = 12'h84D;
            14'd 8490: out = 12'h84D;
            14'd 8491: out = 12'h84E;
            14'd 8492: out = 12'h84E;
            14'd 8493: out = 12'h84E;
            14'd 8494: out = 12'h84E;
            14'd 8495: out = 12'h84F;
            14'd 8496: out = 12'h84F;
            14'd 8497: out = 12'h84F;
            14'd 8498: out = 12'h84F;
            14'd 8499: out = 12'h850;
            14'd 8500: out = 12'h850;
            14'd 8501: out = 12'h850;
            14'd 8502: out = 12'h851;
            14'd 8503: out = 12'h851;
            14'd 8504: out = 12'h851;
            14'd 8505: out = 12'h851;
            14'd 8506: out = 12'h852;
            14'd 8507: out = 12'h852;
            14'd 8508: out = 12'h852;
            14'd 8509: out = 12'h852;
            14'd 8510: out = 12'h853;
            14'd 8511: out = 12'h853;
            14'd 8512: out = 12'h853;
            14'd 8513: out = 12'h854;
            14'd 8514: out = 12'h854;
            14'd 8515: out = 12'h854;
            14'd 8516: out = 12'h854;
            14'd 8517: out = 12'h855;
            14'd 8518: out = 12'h855;
            14'd 8519: out = 12'h855;
            14'd 8520: out = 12'h855;
            14'd 8521: out = 12'h856;
            14'd 8522: out = 12'h856;
            14'd 8523: out = 12'h856;
            14'd 8524: out = 12'h857;
            14'd 8525: out = 12'h857;
            14'd 8526: out = 12'h857;
            14'd 8527: out = 12'h857;
            14'd 8528: out = 12'h858;
            14'd 8529: out = 12'h858;
            14'd 8530: out = 12'h858;
            14'd 8531: out = 12'h858;
            14'd 8532: out = 12'h859;
            14'd 8533: out = 12'h859;
            14'd 8534: out = 12'h859;
            14'd 8535: out = 12'h859;
            14'd 8536: out = 12'h85A;
            14'd 8537: out = 12'h85A;
            14'd 8538: out = 12'h85A;
            14'd 8539: out = 12'h85B;
            14'd 8540: out = 12'h85B;
            14'd 8541: out = 12'h85B;
            14'd 8542: out = 12'h85B;
            14'd 8543: out = 12'h85C;
            14'd 8544: out = 12'h85C;
            14'd 8545: out = 12'h85C;
            14'd 8546: out = 12'h85C;
            14'd 8547: out = 12'h85D;
            14'd 8548: out = 12'h85D;
            14'd 8549: out = 12'h85D;
            14'd 8550: out = 12'h85E;
            14'd 8551: out = 12'h85E;
            14'd 8552: out = 12'h85E;
            14'd 8553: out = 12'h85E;
            14'd 8554: out = 12'h85F;
            14'd 8555: out = 12'h85F;
            14'd 8556: out = 12'h85F;
            14'd 8557: out = 12'h860;
            14'd 8558: out = 12'h860;
            14'd 8559: out = 12'h860;
            14'd 8560: out = 12'h860;
            14'd 8561: out = 12'h861;
            14'd 8562: out = 12'h861;
            14'd 8563: out = 12'h861;
            14'd 8564: out = 12'h861;
            14'd 8565: out = 12'h862;
            14'd 8566: out = 12'h862;
            14'd 8567: out = 12'h862;
            14'd 8568: out = 12'h863;
            14'd 8569: out = 12'h863;
            14'd 8570: out = 12'h863;
            14'd 8571: out = 12'h863;
            14'd 8572: out = 12'h864;
            14'd 8573: out = 12'h864;
            14'd 8574: out = 12'h864;
            14'd 8575: out = 12'h864;
            14'd 8576: out = 12'h865;
            14'd 8577: out = 12'h865;
            14'd 8578: out = 12'h865;
            14'd 8579: out = 12'h866;
            14'd 8580: out = 12'h866;
            14'd 8581: out = 12'h866;
            14'd 8582: out = 12'h866;
            14'd 8583: out = 12'h867;
            14'd 8584: out = 12'h867;
            14'd 8585: out = 12'h867;
            14'd 8586: out = 12'h867;
            14'd 8587: out = 12'h868;
            14'd 8588: out = 12'h868;
            14'd 8589: out = 12'h868;
            14'd 8590: out = 12'h869;
            14'd 8591: out = 12'h869;
            14'd 8592: out = 12'h869;
            14'd 8593: out = 12'h869;
            14'd 8594: out = 12'h86A;
            14'd 8595: out = 12'h86A;
            14'd 8596: out = 12'h86A;
            14'd 8597: out = 12'h86B;
            14'd 8598: out = 12'h86B;
            14'd 8599: out = 12'h86B;
            14'd 8600: out = 12'h86B;
            14'd 8601: out = 12'h86C;
            14'd 8602: out = 12'h86C;
            14'd 8603: out = 12'h86C;
            14'd 8604: out = 12'h86C;
            14'd 8605: out = 12'h86D;
            14'd 8606: out = 12'h86D;
            14'd 8607: out = 12'h86D;
            14'd 8608: out = 12'h86E;
            14'd 8609: out = 12'h86E;
            14'd 8610: out = 12'h86E;
            14'd 8611: out = 12'h86E;
            14'd 8612: out = 12'h86F;
            14'd 8613: out = 12'h86F;
            14'd 8614: out = 12'h86F;
            14'd 8615: out = 12'h870;
            14'd 8616: out = 12'h870;
            14'd 8617: out = 12'h870;
            14'd 8618: out = 12'h870;
            14'd 8619: out = 12'h871;
            14'd 8620: out = 12'h871;
            14'd 8621: out = 12'h871;
            14'd 8622: out = 12'h871;
            14'd 8623: out = 12'h872;
            14'd 8624: out = 12'h872;
            14'd 8625: out = 12'h872;
            14'd 8626: out = 12'h873;
            14'd 8627: out = 12'h873;
            14'd 8628: out = 12'h873;
            14'd 8629: out = 12'h873;
            14'd 8630: out = 12'h874;
            14'd 8631: out = 12'h874;
            14'd 8632: out = 12'h874;
            14'd 8633: out = 12'h875;
            14'd 8634: out = 12'h875;
            14'd 8635: out = 12'h875;
            14'd 8636: out = 12'h875;
            14'd 8637: out = 12'h876;
            14'd 8638: out = 12'h876;
            14'd 8639: out = 12'h876;
            14'd 8640: out = 12'h876;
            14'd 8641: out = 12'h877;
            14'd 8642: out = 12'h877;
            14'd 8643: out = 12'h877;
            14'd 8644: out = 12'h878;
            14'd 8645: out = 12'h878;
            14'd 8646: out = 12'h878;
            14'd 8647: out = 12'h878;
            14'd 8648: out = 12'h879;
            14'd 8649: out = 12'h879;
            14'd 8650: out = 12'h879;
            14'd 8651: out = 12'h87A;
            14'd 8652: out = 12'h87A;
            14'd 8653: out = 12'h87A;
            14'd 8654: out = 12'h87A;
            14'd 8655: out = 12'h87B;
            14'd 8656: out = 12'h87B;
            14'd 8657: out = 12'h87B;
            14'd 8658: out = 12'h87C;
            14'd 8659: out = 12'h87C;
            14'd 8660: out = 12'h87C;
            14'd 8661: out = 12'h87C;
            14'd 8662: out = 12'h87D;
            14'd 8663: out = 12'h87D;
            14'd 8664: out = 12'h87D;
            14'd 8665: out = 12'h87D;
            14'd 8666: out = 12'h87E;
            14'd 8667: out = 12'h87E;
            14'd 8668: out = 12'h87E;
            14'd 8669: out = 12'h87F;
            14'd 8670: out = 12'h87F;
            14'd 8671: out = 12'h87F;
            14'd 8672: out = 12'h87F;
            14'd 8673: out = 12'h880;
            14'd 8674: out = 12'h880;
            14'd 8675: out = 12'h880;
            14'd 8676: out = 12'h881;
            14'd 8677: out = 12'h881;
            14'd 8678: out = 12'h881;
            14'd 8679: out = 12'h881;
            14'd 8680: out = 12'h882;
            14'd 8681: out = 12'h882;
            14'd 8682: out = 12'h882;
            14'd 8683: out = 12'h883;
            14'd 8684: out = 12'h883;
            14'd 8685: out = 12'h883;
            14'd 8686: out = 12'h883;
            14'd 8687: out = 12'h884;
            14'd 8688: out = 12'h884;
            14'd 8689: out = 12'h884;
            14'd 8690: out = 12'h885;
            14'd 8691: out = 12'h885;
            14'd 8692: out = 12'h885;
            14'd 8693: out = 12'h885;
            14'd 8694: out = 12'h886;
            14'd 8695: out = 12'h886;
            14'd 8696: out = 12'h886;
            14'd 8697: out = 12'h887;
            14'd 8698: out = 12'h887;
            14'd 8699: out = 12'h887;
            14'd 8700: out = 12'h887;
            14'd 8701: out = 12'h888;
            14'd 8702: out = 12'h888;
            14'd 8703: out = 12'h888;
            14'd 8704: out = 12'h889;
            14'd 8705: out = 12'h889;
            14'd 8706: out = 12'h889;
            14'd 8707: out = 12'h889;
            14'd 8708: out = 12'h88A;
            14'd 8709: out = 12'h88A;
            14'd 8710: out = 12'h88A;
            14'd 8711: out = 12'h88B;
            14'd 8712: out = 12'h88B;
            14'd 8713: out = 12'h88B;
            14'd 8714: out = 12'h88B;
            14'd 8715: out = 12'h88C;
            14'd 8716: out = 12'h88C;
            14'd 8717: out = 12'h88C;
            14'd 8718: out = 12'h88D;
            14'd 8719: out = 12'h88D;
            14'd 8720: out = 12'h88D;
            14'd 8721: out = 12'h88D;
            14'd 8722: out = 12'h88E;
            14'd 8723: out = 12'h88E;
            14'd 8724: out = 12'h88E;
            14'd 8725: out = 12'h88F;
            14'd 8726: out = 12'h88F;
            14'd 8727: out = 12'h88F;
            14'd 8728: out = 12'h88F;
            14'd 8729: out = 12'h890;
            14'd 8730: out = 12'h890;
            14'd 8731: out = 12'h890;
            14'd 8732: out = 12'h891;
            14'd 8733: out = 12'h891;
            14'd 8734: out = 12'h891;
            14'd 8735: out = 12'h891;
            14'd 8736: out = 12'h892;
            14'd 8737: out = 12'h892;
            14'd 8738: out = 12'h892;
            14'd 8739: out = 12'h893;
            14'd 8740: out = 12'h893;
            14'd 8741: out = 12'h893;
            14'd 8742: out = 12'h893;
            14'd 8743: out = 12'h894;
            14'd 8744: out = 12'h894;
            14'd 8745: out = 12'h894;
            14'd 8746: out = 12'h895;
            14'd 8747: out = 12'h895;
            14'd 8748: out = 12'h895;
            14'd 8749: out = 12'h895;
            14'd 8750: out = 12'h896;
            14'd 8751: out = 12'h896;
            14'd 8752: out = 12'h896;
            14'd 8753: out = 12'h897;
            14'd 8754: out = 12'h897;
            14'd 8755: out = 12'h897;
            14'd 8756: out = 12'h897;
            14'd 8757: out = 12'h898;
            14'd 8758: out = 12'h898;
            14'd 8759: out = 12'h898;
            14'd 8760: out = 12'h899;
            14'd 8761: out = 12'h899;
            14'd 8762: out = 12'h899;
            14'd 8763: out = 12'h899;
            14'd 8764: out = 12'h89A;
            14'd 8765: out = 12'h89A;
            14'd 8766: out = 12'h89A;
            14'd 8767: out = 12'h89B;
            14'd 8768: out = 12'h89B;
            14'd 8769: out = 12'h89B;
            14'd 8770: out = 12'h89B;
            14'd 8771: out = 12'h89C;
            14'd 8772: out = 12'h89C;
            14'd 8773: out = 12'h89C;
            14'd 8774: out = 12'h89D;
            14'd 8775: out = 12'h89D;
            14'd 8776: out = 12'h89D;
            14'd 8777: out = 12'h89D;
            14'd 8778: out = 12'h89E;
            14'd 8779: out = 12'h89E;
            14'd 8780: out = 12'h89E;
            14'd 8781: out = 12'h89F;
            14'd 8782: out = 12'h89F;
            14'd 8783: out = 12'h89F;
            14'd 8784: out = 12'h8A0;
            14'd 8785: out = 12'h8A0;
            14'd 8786: out = 12'h8A0;
            14'd 8787: out = 12'h8A0;
            14'd 8788: out = 12'h8A1;
            14'd 8789: out = 12'h8A1;
            14'd 8790: out = 12'h8A1;
            14'd 8791: out = 12'h8A2;
            14'd 8792: out = 12'h8A2;
            14'd 8793: out = 12'h8A2;
            14'd 8794: out = 12'h8A2;
            14'd 8795: out = 12'h8A3;
            14'd 8796: out = 12'h8A3;
            14'd 8797: out = 12'h8A3;
            14'd 8798: out = 12'h8A4;
            14'd 8799: out = 12'h8A4;
            14'd 8800: out = 12'h8A4;
            14'd 8801: out = 12'h8A4;
            14'd 8802: out = 12'h8A5;
            14'd 8803: out = 12'h8A5;
            14'd 8804: out = 12'h8A5;
            14'd 8805: out = 12'h8A6;
            14'd 8806: out = 12'h8A6;
            14'd 8807: out = 12'h8A6;
            14'd 8808: out = 12'h8A7;
            14'd 8809: out = 12'h8A7;
            14'd 8810: out = 12'h8A7;
            14'd 8811: out = 12'h8A7;
            14'd 8812: out = 12'h8A8;
            14'd 8813: out = 12'h8A8;
            14'd 8814: out = 12'h8A8;
            14'd 8815: out = 12'h8A9;
            14'd 8816: out = 12'h8A9;
            14'd 8817: out = 12'h8A9;
            14'd 8818: out = 12'h8A9;
            14'd 8819: out = 12'h8AA;
            14'd 8820: out = 12'h8AA;
            14'd 8821: out = 12'h8AA;
            14'd 8822: out = 12'h8AB;
            14'd 8823: out = 12'h8AB;
            14'd 8824: out = 12'h8AB;
            14'd 8825: out = 12'h8AC;
            14'd 8826: out = 12'h8AC;
            14'd 8827: out = 12'h8AC;
            14'd 8828: out = 12'h8AC;
            14'd 8829: out = 12'h8AD;
            14'd 8830: out = 12'h8AD;
            14'd 8831: out = 12'h8AD;
            14'd 8832: out = 12'h8AE;
            14'd 8833: out = 12'h8AE;
            14'd 8834: out = 12'h8AE;
            14'd 8835: out = 12'h8AE;
            14'd 8836: out = 12'h8AF;
            14'd 8837: out = 12'h8AF;
            14'd 8838: out = 12'h8AF;
            14'd 8839: out = 12'h8B0;
            14'd 8840: out = 12'h8B0;
            14'd 8841: out = 12'h8B0;
            14'd 8842: out = 12'h8B1;
            14'd 8843: out = 12'h8B1;
            14'd 8844: out = 12'h8B1;
            14'd 8845: out = 12'h8B1;
            14'd 8846: out = 12'h8B2;
            14'd 8847: out = 12'h8B2;
            14'd 8848: out = 12'h8B2;
            14'd 8849: out = 12'h8B3;
            14'd 8850: out = 12'h8B3;
            14'd 8851: out = 12'h8B3;
            14'd 8852: out = 12'h8B3;
            14'd 8853: out = 12'h8B4;
            14'd 8854: out = 12'h8B4;
            14'd 8855: out = 12'h8B4;
            14'd 8856: out = 12'h8B5;
            14'd 8857: out = 12'h8B5;
            14'd 8858: out = 12'h8B5;
            14'd 8859: out = 12'h8B6;
            14'd 8860: out = 12'h8B6;
            14'd 8861: out = 12'h8B6;
            14'd 8862: out = 12'h8B6;
            14'd 8863: out = 12'h8B7;
            14'd 8864: out = 12'h8B7;
            14'd 8865: out = 12'h8B7;
            14'd 8866: out = 12'h8B8;
            14'd 8867: out = 12'h8B8;
            14'd 8868: out = 12'h8B8;
            14'd 8869: out = 12'h8B8;
            14'd 8870: out = 12'h8B9;
            14'd 8871: out = 12'h8B9;
            14'd 8872: out = 12'h8B9;
            14'd 8873: out = 12'h8BA;
            14'd 8874: out = 12'h8BA;
            14'd 8875: out = 12'h8BA;
            14'd 8876: out = 12'h8BB;
            14'd 8877: out = 12'h8BB;
            14'd 8878: out = 12'h8BB;
            14'd 8879: out = 12'h8BB;
            14'd 8880: out = 12'h8BC;
            14'd 8881: out = 12'h8BC;
            14'd 8882: out = 12'h8BC;
            14'd 8883: out = 12'h8BD;
            14'd 8884: out = 12'h8BD;
            14'd 8885: out = 12'h8BD;
            14'd 8886: out = 12'h8BE;
            14'd 8887: out = 12'h8BE;
            14'd 8888: out = 12'h8BE;
            14'd 8889: out = 12'h8BE;
            14'd 8890: out = 12'h8BF;
            14'd 8891: out = 12'h8BF;
            14'd 8892: out = 12'h8BF;
            14'd 8893: out = 12'h8C0;
            14'd 8894: out = 12'h8C0;
            14'd 8895: out = 12'h8C0;
            14'd 8896: out = 12'h8C1;
            14'd 8897: out = 12'h8C1;
            14'd 8898: out = 12'h8C1;
            14'd 8899: out = 12'h8C1;
            14'd 8900: out = 12'h8C2;
            14'd 8901: out = 12'h8C2;
            14'd 8902: out = 12'h8C2;
            14'd 8903: out = 12'h8C3;
            14'd 8904: out = 12'h8C3;
            14'd 8905: out = 12'h8C3;
            14'd 8906: out = 12'h8C4;
            14'd 8907: out = 12'h8C4;
            14'd 8908: out = 12'h8C4;
            14'd 8909: out = 12'h8C4;
            14'd 8910: out = 12'h8C5;
            14'd 8911: out = 12'h8C5;
            14'd 8912: out = 12'h8C5;
            14'd 8913: out = 12'h8C6;
            14'd 8914: out = 12'h8C6;
            14'd 8915: out = 12'h8C6;
            14'd 8916: out = 12'h8C7;
            14'd 8917: out = 12'h8C7;
            14'd 8918: out = 12'h8C7;
            14'd 8919: out = 12'h8C7;
            14'd 8920: out = 12'h8C8;
            14'd 8921: out = 12'h8C8;
            14'd 8922: out = 12'h8C8;
            14'd 8923: out = 12'h8C9;
            14'd 8924: out = 12'h8C9;
            14'd 8925: out = 12'h8C9;
            14'd 8926: out = 12'h8CA;
            14'd 8927: out = 12'h8CA;
            14'd 8928: out = 12'h8CA;
            14'd 8929: out = 12'h8CA;
            14'd 8930: out = 12'h8CB;
            14'd 8931: out = 12'h8CB;
            14'd 8932: out = 12'h8CB;
            14'd 8933: out = 12'h8CC;
            14'd 8934: out = 12'h8CC;
            14'd 8935: out = 12'h8CC;
            14'd 8936: out = 12'h8CD;
            14'd 8937: out = 12'h8CD;
            14'd 8938: out = 12'h8CD;
            14'd 8939: out = 12'h8CD;
            14'd 8940: out = 12'h8CE;
            14'd 8941: out = 12'h8CE;
            14'd 8942: out = 12'h8CE;
            14'd 8943: out = 12'h8CF;
            14'd 8944: out = 12'h8CF;
            14'd 8945: out = 12'h8CF;
            14'd 8946: out = 12'h8D0;
            14'd 8947: out = 12'h8D0;
            14'd 8948: out = 12'h8D0;
            14'd 8949: out = 12'h8D1;
            14'd 8950: out = 12'h8D1;
            14'd 8951: out = 12'h8D1;
            14'd 8952: out = 12'h8D1;
            14'd 8953: out = 12'h8D2;
            14'd 8954: out = 12'h8D2;
            14'd 8955: out = 12'h8D2;
            14'd 8956: out = 12'h8D3;
            14'd 8957: out = 12'h8D3;
            14'd 8958: out = 12'h8D3;
            14'd 8959: out = 12'h8D4;
            14'd 8960: out = 12'h8D4;
            14'd 8961: out = 12'h8D4;
            14'd 8962: out = 12'h8D4;
            14'd 8963: out = 12'h8D5;
            14'd 8964: out = 12'h8D5;
            14'd 8965: out = 12'h8D5;
            14'd 8966: out = 12'h8D6;
            14'd 8967: out = 12'h8D6;
            14'd 8968: out = 12'h8D6;
            14'd 8969: out = 12'h8D7;
            14'd 8970: out = 12'h8D7;
            14'd 8971: out = 12'h8D7;
            14'd 8972: out = 12'h8D8;
            14'd 8973: out = 12'h8D8;
            14'd 8974: out = 12'h8D8;
            14'd 8975: out = 12'h8D8;
            14'd 8976: out = 12'h8D9;
            14'd 8977: out = 12'h8D9;
            14'd 8978: out = 12'h8D9;
            14'd 8979: out = 12'h8DA;
            14'd 8980: out = 12'h8DA;
            14'd 8981: out = 12'h8DA;
            14'd 8982: out = 12'h8DB;
            14'd 8983: out = 12'h8DB;
            14'd 8984: out = 12'h8DB;
            14'd 8985: out = 12'h8DB;
            14'd 8986: out = 12'h8DC;
            14'd 8987: out = 12'h8DC;
            14'd 8988: out = 12'h8DC;
            14'd 8989: out = 12'h8DD;
            14'd 8990: out = 12'h8DD;
            14'd 8991: out = 12'h8DD;
            14'd 8992: out = 12'h8DE;
            14'd 8993: out = 12'h8DE;
            14'd 8994: out = 12'h8DE;
            14'd 8995: out = 12'h8DF;
            14'd 8996: out = 12'h8DF;
            14'd 8997: out = 12'h8DF;
            14'd 8998: out = 12'h8DF;
            14'd 8999: out = 12'h8E0;
            14'd 9000: out = 12'h8E0;
            14'd 9001: out = 12'h8E0;
            14'd 9002: out = 12'h8E1;
            14'd 9003: out = 12'h8E1;
            14'd 9004: out = 12'h8E1;
            14'd 9005: out = 12'h8E2;
            14'd 9006: out = 12'h8E2;
            14'd 9007: out = 12'h8E2;
            14'd 9008: out = 12'h8E3;
            14'd 9009: out = 12'h8E3;
            14'd 9010: out = 12'h8E3;
            14'd 9011: out = 12'h8E3;
            14'd 9012: out = 12'h8E4;
            14'd 9013: out = 12'h8E4;
            14'd 9014: out = 12'h8E4;
            14'd 9015: out = 12'h8E5;
            14'd 9016: out = 12'h8E5;
            14'd 9017: out = 12'h8E5;
            14'd 9018: out = 12'h8E6;
            14'd 9019: out = 12'h8E6;
            14'd 9020: out = 12'h8E6;
            14'd 9021: out = 12'h8E7;
            14'd 9022: out = 12'h8E7;
            14'd 9023: out = 12'h8E7;
            14'd 9024: out = 12'h8E8;
            14'd 9025: out = 12'h8E8;
            14'd 9026: out = 12'h8E8;
            14'd 9027: out = 12'h8E8;
            14'd 9028: out = 12'h8E9;
            14'd 9029: out = 12'h8E9;
            14'd 9030: out = 12'h8E9;
            14'd 9031: out = 12'h8EA;
            14'd 9032: out = 12'h8EA;
            14'd 9033: out = 12'h8EA;
            14'd 9034: out = 12'h8EB;
            14'd 9035: out = 12'h8EB;
            14'd 9036: out = 12'h8EB;
            14'd 9037: out = 12'h8EC;
            14'd 9038: out = 12'h8EC;
            14'd 9039: out = 12'h8EC;
            14'd 9040: out = 12'h8EC;
            14'd 9041: out = 12'h8ED;
            14'd 9042: out = 12'h8ED;
            14'd 9043: out = 12'h8ED;
            14'd 9044: out = 12'h8EE;
            14'd 9045: out = 12'h8EE;
            14'd 9046: out = 12'h8EE;
            14'd 9047: out = 12'h8EF;
            14'd 9048: out = 12'h8EF;
            14'd 9049: out = 12'h8EF;
            14'd 9050: out = 12'h8F0;
            14'd 9051: out = 12'h8F0;
            14'd 9052: out = 12'h8F0;
            14'd 9053: out = 12'h8F1;
            14'd 9054: out = 12'h8F1;
            14'd 9055: out = 12'h8F1;
            14'd 9056: out = 12'h8F1;
            14'd 9057: out = 12'h8F2;
            14'd 9058: out = 12'h8F2;
            14'd 9059: out = 12'h8F2;
            14'd 9060: out = 12'h8F3;
            14'd 9061: out = 12'h8F3;
            14'd 9062: out = 12'h8F3;
            14'd 9063: out = 12'h8F4;
            14'd 9064: out = 12'h8F4;
            14'd 9065: out = 12'h8F4;
            14'd 9066: out = 12'h8F5;
            14'd 9067: out = 12'h8F5;
            14'd 9068: out = 12'h8F5;
            14'd 9069: out = 12'h8F6;
            14'd 9070: out = 12'h8F6;
            14'd 9071: out = 12'h8F6;
            14'd 9072: out = 12'h8F6;
            14'd 9073: out = 12'h8F7;
            14'd 9074: out = 12'h8F7;
            14'd 9075: out = 12'h8F7;
            14'd 9076: out = 12'h8F8;
            14'd 9077: out = 12'h8F8;
            14'd 9078: out = 12'h8F8;
            14'd 9079: out = 12'h8F9;
            14'd 9080: out = 12'h8F9;
            14'd 9081: out = 12'h8F9;
            14'd 9082: out = 12'h8FA;
            14'd 9083: out = 12'h8FA;
            14'd 9084: out = 12'h8FA;
            14'd 9085: out = 12'h8FB;
            14'd 9086: out = 12'h8FB;
            14'd 9087: out = 12'h8FB;
            14'd 9088: out = 12'h8FC;
            14'd 9089: out = 12'h8FC;
            14'd 9090: out = 12'h8FC;
            14'd 9091: out = 12'h8FC;
            14'd 9092: out = 12'h8FD;
            14'd 9093: out = 12'h8FD;
            14'd 9094: out = 12'h8FD;
            14'd 9095: out = 12'h8FE;
            14'd 9096: out = 12'h8FE;
            14'd 9097: out = 12'h8FE;
            14'd 9098: out = 12'h8FF;
            14'd 9099: out = 12'h8FF;
            14'd 9100: out = 12'h8FF;
            14'd 9101: out = 12'h900;
            14'd 9102: out = 12'h900;
            14'd 9103: out = 12'h900;
            14'd 9104: out = 12'h901;
            14'd 9105: out = 12'h901;
            14'd 9106: out = 12'h901;
            14'd 9107: out = 12'h902;
            14'd 9108: out = 12'h902;
            14'd 9109: out = 12'h902;
            14'd 9110: out = 12'h902;
            14'd 9111: out = 12'h903;
            14'd 9112: out = 12'h903;
            14'd 9113: out = 12'h903;
            14'd 9114: out = 12'h904;
            14'd 9115: out = 12'h904;
            14'd 9116: out = 12'h904;
            14'd 9117: out = 12'h905;
            14'd 9118: out = 12'h905;
            14'd 9119: out = 12'h905;
            14'd 9120: out = 12'h906;
            14'd 9121: out = 12'h906;
            14'd 9122: out = 12'h906;
            14'd 9123: out = 12'h907;
            14'd 9124: out = 12'h907;
            14'd 9125: out = 12'h907;
            14'd 9126: out = 12'h908;
            14'd 9127: out = 12'h908;
            14'd 9128: out = 12'h908;
            14'd 9129: out = 12'h909;
            14'd 9130: out = 12'h909;
            14'd 9131: out = 12'h909;
            14'd 9132: out = 12'h909;
            14'd 9133: out = 12'h90A;
            14'd 9134: out = 12'h90A;
            14'd 9135: out = 12'h90A;
            14'd 9136: out = 12'h90B;
            14'd 9137: out = 12'h90B;
            14'd 9138: out = 12'h90B;
            14'd 9139: out = 12'h90C;
            14'd 9140: out = 12'h90C;
            14'd 9141: out = 12'h90C;
            14'd 9142: out = 12'h90D;
            14'd 9143: out = 12'h90D;
            14'd 9144: out = 12'h90D;
            14'd 9145: out = 12'h90E;
            14'd 9146: out = 12'h90E;
            14'd 9147: out = 12'h90E;
            14'd 9148: out = 12'h90F;
            14'd 9149: out = 12'h90F;
            14'd 9150: out = 12'h90F;
            14'd 9151: out = 12'h910;
            14'd 9152: out = 12'h910;
            14'd 9153: out = 12'h910;
            14'd 9154: out = 12'h911;
            14'd 9155: out = 12'h911;
            14'd 9156: out = 12'h911;
            14'd 9157: out = 12'h911;
            14'd 9158: out = 12'h912;
            14'd 9159: out = 12'h912;
            14'd 9160: out = 12'h912;
            14'd 9161: out = 12'h913;
            14'd 9162: out = 12'h913;
            14'd 9163: out = 12'h913;
            14'd 9164: out = 12'h914;
            14'd 9165: out = 12'h914;
            14'd 9166: out = 12'h914;
            14'd 9167: out = 12'h915;
            14'd 9168: out = 12'h915;
            14'd 9169: out = 12'h915;
            14'd 9170: out = 12'h916;
            14'd 9171: out = 12'h916;
            14'd 9172: out = 12'h916;
            14'd 9173: out = 12'h917;
            14'd 9174: out = 12'h917;
            14'd 9175: out = 12'h917;
            14'd 9176: out = 12'h918;
            14'd 9177: out = 12'h918;
            14'd 9178: out = 12'h918;
            14'd 9179: out = 12'h919;
            14'd 9180: out = 12'h919;
            14'd 9181: out = 12'h919;
            14'd 9182: out = 12'h91A;
            14'd 9183: out = 12'h91A;
            14'd 9184: out = 12'h91A;
            14'd 9185: out = 12'h91A;
            14'd 9186: out = 12'h91B;
            14'd 9187: out = 12'h91B;
            14'd 9188: out = 12'h91B;
            14'd 9189: out = 12'h91C;
            14'd 9190: out = 12'h91C;
            14'd 9191: out = 12'h91C;
            14'd 9192: out = 12'h91D;
            14'd 9193: out = 12'h91D;
            14'd 9194: out = 12'h91D;
            14'd 9195: out = 12'h91E;
            14'd 9196: out = 12'h91E;
            14'd 9197: out = 12'h91E;
            14'd 9198: out = 12'h91F;
            14'd 9199: out = 12'h91F;
            14'd 9200: out = 12'h91F;
            14'd 9201: out = 12'h920;
            14'd 9202: out = 12'h920;
            14'd 9203: out = 12'h920;
            14'd 9204: out = 12'h921;
            14'd 9205: out = 12'h921;
            14'd 9206: out = 12'h921;
            14'd 9207: out = 12'h922;
            14'd 9208: out = 12'h922;
            14'd 9209: out = 12'h922;
            14'd 9210: out = 12'h923;
            14'd 9211: out = 12'h923;
            14'd 9212: out = 12'h923;
            14'd 9213: out = 12'h924;
            14'd 9214: out = 12'h924;
            14'd 9215: out = 12'h924;
            14'd 9216: out = 12'h925;
            14'd 9217: out = 12'h925;
            14'd 9218: out = 12'h925;
            14'd 9219: out = 12'h926;
            14'd 9220: out = 12'h926;
            14'd 9221: out = 12'h926;
            14'd 9222: out = 12'h927;
            14'd 9223: out = 12'h927;
            14'd 9224: out = 12'h927;
            14'd 9225: out = 12'h928;
            14'd 9226: out = 12'h928;
            14'd 9227: out = 12'h928;
            14'd 9228: out = 12'h928;
            14'd 9229: out = 12'h929;
            14'd 9230: out = 12'h929;
            14'd 9231: out = 12'h929;
            14'd 9232: out = 12'h92A;
            14'd 9233: out = 12'h92A;
            14'd 9234: out = 12'h92A;
            14'd 9235: out = 12'h92B;
            14'd 9236: out = 12'h92B;
            14'd 9237: out = 12'h92B;
            14'd 9238: out = 12'h92C;
            14'd 9239: out = 12'h92C;
            14'd 9240: out = 12'h92C;
            14'd 9241: out = 12'h92D;
            14'd 9242: out = 12'h92D;
            14'd 9243: out = 12'h92D;
            14'd 9244: out = 12'h92E;
            14'd 9245: out = 12'h92E;
            14'd 9246: out = 12'h92E;
            14'd 9247: out = 12'h92F;
            14'd 9248: out = 12'h92F;
            14'd 9249: out = 12'h92F;
            14'd 9250: out = 12'h930;
            14'd 9251: out = 12'h930;
            14'd 9252: out = 12'h930;
            14'd 9253: out = 12'h931;
            14'd 9254: out = 12'h931;
            14'd 9255: out = 12'h931;
            14'd 9256: out = 12'h932;
            14'd 9257: out = 12'h932;
            14'd 9258: out = 12'h932;
            14'd 9259: out = 12'h933;
            14'd 9260: out = 12'h933;
            14'd 9261: out = 12'h933;
            14'd 9262: out = 12'h934;
            14'd 9263: out = 12'h934;
            14'd 9264: out = 12'h934;
            14'd 9265: out = 12'h935;
            14'd 9266: out = 12'h935;
            14'd 9267: out = 12'h935;
            14'd 9268: out = 12'h936;
            14'd 9269: out = 12'h936;
            14'd 9270: out = 12'h936;
            14'd 9271: out = 12'h937;
            14'd 9272: out = 12'h937;
            14'd 9273: out = 12'h937;
            14'd 9274: out = 12'h938;
            14'd 9275: out = 12'h938;
            14'd 9276: out = 12'h938;
            14'd 9277: out = 12'h939;
            14'd 9278: out = 12'h939;
            14'd 9279: out = 12'h939;
            14'd 9280: out = 12'h93A;
            14'd 9281: out = 12'h93A;
            14'd 9282: out = 12'h93A;
            14'd 9283: out = 12'h93B;
            14'd 9284: out = 12'h93B;
            14'd 9285: out = 12'h93B;
            14'd 9286: out = 12'h93C;
            14'd 9287: out = 12'h93C;
            14'd 9288: out = 12'h93C;
            14'd 9289: out = 12'h93D;
            14'd 9290: out = 12'h93D;
            14'd 9291: out = 12'h93D;
            14'd 9292: out = 12'h93E;
            14'd 9293: out = 12'h93E;
            14'd 9294: out = 12'h93E;
            14'd 9295: out = 12'h93F;
            14'd 9296: out = 12'h93F;
            14'd 9297: out = 12'h93F;
            14'd 9298: out = 12'h940;
            14'd 9299: out = 12'h940;
            14'd 9300: out = 12'h940;
            14'd 9301: out = 12'h941;
            14'd 9302: out = 12'h941;
            14'd 9303: out = 12'h941;
            14'd 9304: out = 12'h942;
            14'd 9305: out = 12'h942;
            14'd 9306: out = 12'h942;
            14'd 9307: out = 12'h943;
            14'd 9308: out = 12'h943;
            14'd 9309: out = 12'h943;
            14'd 9310: out = 12'h944;
            14'd 9311: out = 12'h944;
            14'd 9312: out = 12'h944;
            14'd 9313: out = 12'h945;
            14'd 9314: out = 12'h945;
            14'd 9315: out = 12'h945;
            14'd 9316: out = 12'h946;
            14'd 9317: out = 12'h946;
            14'd 9318: out = 12'h946;
            14'd 9319: out = 12'h947;
            14'd 9320: out = 12'h947;
            14'd 9321: out = 12'h947;
            14'd 9322: out = 12'h948;
            14'd 9323: out = 12'h948;
            14'd 9324: out = 12'h948;
            14'd 9325: out = 12'h949;
            14'd 9326: out = 12'h949;
            14'd 9327: out = 12'h949;
            14'd 9328: out = 12'h94A;
            14'd 9329: out = 12'h94A;
            14'd 9330: out = 12'h94A;
            14'd 9331: out = 12'h94B;
            14'd 9332: out = 12'h94B;
            14'd 9333: out = 12'h94B;
            14'd 9334: out = 12'h94C;
            14'd 9335: out = 12'h94C;
            14'd 9336: out = 12'h94C;
            14'd 9337: out = 12'h94D;
            14'd 9338: out = 12'h94D;
            14'd 9339: out = 12'h94D;
            14'd 9340: out = 12'h94E;
            14'd 9341: out = 12'h94E;
            14'd 9342: out = 12'h94E;
            14'd 9343: out = 12'h94F;
            14'd 9344: out = 12'h94F;
            14'd 9345: out = 12'h94F;
            14'd 9346: out = 12'h950;
            14'd 9347: out = 12'h950;
            14'd 9348: out = 12'h950;
            14'd 9349: out = 12'h951;
            14'd 9350: out = 12'h951;
            14'd 9351: out = 12'h951;
            14'd 9352: out = 12'h952;
            14'd 9353: out = 12'h952;
            14'd 9354: out = 12'h953;
            14'd 9355: out = 12'h953;
            14'd 9356: out = 12'h953;
            14'd 9357: out = 12'h954;
            14'd 9358: out = 12'h954;
            14'd 9359: out = 12'h954;
            14'd 9360: out = 12'h955;
            14'd 9361: out = 12'h955;
            14'd 9362: out = 12'h955;
            14'd 9363: out = 12'h956;
            14'd 9364: out = 12'h956;
            14'd 9365: out = 12'h956;
            14'd 9366: out = 12'h957;
            14'd 9367: out = 12'h957;
            14'd 9368: out = 12'h957;
            14'd 9369: out = 12'h958;
            14'd 9370: out = 12'h958;
            14'd 9371: out = 12'h958;
            14'd 9372: out = 12'h959;
            14'd 9373: out = 12'h959;
            14'd 9374: out = 12'h959;
            14'd 9375: out = 12'h95A;
            14'd 9376: out = 12'h95A;
            14'd 9377: out = 12'h95A;
            14'd 9378: out = 12'h95B;
            14'd 9379: out = 12'h95B;
            14'd 9380: out = 12'h95B;
            14'd 9381: out = 12'h95C;
            14'd 9382: out = 12'h95C;
            14'd 9383: out = 12'h95C;
            14'd 9384: out = 12'h95D;
            14'd 9385: out = 12'h95D;
            14'd 9386: out = 12'h95D;
            14'd 9387: out = 12'h95E;
            14'd 9388: out = 12'h95E;
            14'd 9389: out = 12'h95E;
            14'd 9390: out = 12'h95F;
            14'd 9391: out = 12'h95F;
            14'd 9392: out = 12'h95F;
            14'd 9393: out = 12'h960;
            14'd 9394: out = 12'h960;
            14'd 9395: out = 12'h961;
            14'd 9396: out = 12'h961;
            14'd 9397: out = 12'h961;
            14'd 9398: out = 12'h962;
            14'd 9399: out = 12'h962;
            14'd 9400: out = 12'h962;
            14'd 9401: out = 12'h963;
            14'd 9402: out = 12'h963;
            14'd 9403: out = 12'h963;
            14'd 9404: out = 12'h964;
            14'd 9405: out = 12'h964;
            14'd 9406: out = 12'h964;
            14'd 9407: out = 12'h965;
            14'd 9408: out = 12'h965;
            14'd 9409: out = 12'h965;
            14'd 9410: out = 12'h966;
            14'd 9411: out = 12'h966;
            14'd 9412: out = 12'h966;
            14'd 9413: out = 12'h967;
            14'd 9414: out = 12'h967;
            14'd 9415: out = 12'h967;
            14'd 9416: out = 12'h968;
            14'd 9417: out = 12'h968;
            14'd 9418: out = 12'h968;
            14'd 9419: out = 12'h969;
            14'd 9420: out = 12'h969;
            14'd 9421: out = 12'h969;
            14'd 9422: out = 12'h96A;
            14'd 9423: out = 12'h96A;
            14'd 9424: out = 12'h96B;
            14'd 9425: out = 12'h96B;
            14'd 9426: out = 12'h96B;
            14'd 9427: out = 12'h96C;
            14'd 9428: out = 12'h96C;
            14'd 9429: out = 12'h96C;
            14'd 9430: out = 12'h96D;
            14'd 9431: out = 12'h96D;
            14'd 9432: out = 12'h96D;
            14'd 9433: out = 12'h96E;
            14'd 9434: out = 12'h96E;
            14'd 9435: out = 12'h96E;
            14'd 9436: out = 12'h96F;
            14'd 9437: out = 12'h96F;
            14'd 9438: out = 12'h96F;
            14'd 9439: out = 12'h970;
            14'd 9440: out = 12'h970;
            14'd 9441: out = 12'h970;
            14'd 9442: out = 12'h971;
            14'd 9443: out = 12'h971;
            14'd 9444: out = 12'h971;
            14'd 9445: out = 12'h972;
            14'd 9446: out = 12'h972;
            14'd 9447: out = 12'h973;
            14'd 9448: out = 12'h973;
            14'd 9449: out = 12'h973;
            14'd 9450: out = 12'h974;
            14'd 9451: out = 12'h974;
            14'd 9452: out = 12'h974;
            14'd 9453: out = 12'h975;
            14'd 9454: out = 12'h975;
            14'd 9455: out = 12'h975;
            14'd 9456: out = 12'h976;
            14'd 9457: out = 12'h976;
            14'd 9458: out = 12'h976;
            14'd 9459: out = 12'h977;
            14'd 9460: out = 12'h977;
            14'd 9461: out = 12'h977;
            14'd 9462: out = 12'h978;
            14'd 9463: out = 12'h978;
            14'd 9464: out = 12'h978;
            14'd 9465: out = 12'h979;
            14'd 9466: out = 12'h979;
            14'd 9467: out = 12'h97A;
            14'd 9468: out = 12'h97A;
            14'd 9469: out = 12'h97A;
            14'd 9470: out = 12'h97B;
            14'd 9471: out = 12'h97B;
            14'd 9472: out = 12'h97B;
            14'd 9473: out = 12'h97C;
            14'd 9474: out = 12'h97C;
            14'd 9475: out = 12'h97C;
            14'd 9476: out = 12'h97D;
            14'd 9477: out = 12'h97D;
            14'd 9478: out = 12'h97D;
            14'd 9479: out = 12'h97E;
            14'd 9480: out = 12'h97E;
            14'd 9481: out = 12'h97E;
            14'd 9482: out = 12'h97F;
            14'd 9483: out = 12'h97F;
            14'd 9484: out = 12'h97F;
            14'd 9485: out = 12'h980;
            14'd 9486: out = 12'h980;
            14'd 9487: out = 12'h981;
            14'd 9488: out = 12'h981;
            14'd 9489: out = 12'h981;
            14'd 9490: out = 12'h982;
            14'd 9491: out = 12'h982;
            14'd 9492: out = 12'h982;
            14'd 9493: out = 12'h983;
            14'd 9494: out = 12'h983;
            14'd 9495: out = 12'h983;
            14'd 9496: out = 12'h984;
            14'd 9497: out = 12'h984;
            14'd 9498: out = 12'h984;
            14'd 9499: out = 12'h985;
            14'd 9500: out = 12'h985;
            14'd 9501: out = 12'h985;
            14'd 9502: out = 12'h986;
            14'd 9503: out = 12'h986;
            14'd 9504: out = 12'h987;
            14'd 9505: out = 12'h987;
            14'd 9506: out = 12'h987;
            14'd 9507: out = 12'h988;
            14'd 9508: out = 12'h988;
            14'd 9509: out = 12'h988;
            14'd 9510: out = 12'h989;
            14'd 9511: out = 12'h989;
            14'd 9512: out = 12'h989;
            14'd 9513: out = 12'h98A;
            14'd 9514: out = 12'h98A;
            14'd 9515: out = 12'h98A;
            14'd 9516: out = 12'h98B;
            14'd 9517: out = 12'h98B;
            14'd 9518: out = 12'h98C;
            14'd 9519: out = 12'h98C;
            14'd 9520: out = 12'h98C;
            14'd 9521: out = 12'h98D;
            14'd 9522: out = 12'h98D;
            14'd 9523: out = 12'h98D;
            14'd 9524: out = 12'h98E;
            14'd 9525: out = 12'h98E;
            14'd 9526: out = 12'h98E;
            14'd 9527: out = 12'h98F;
            14'd 9528: out = 12'h98F;
            14'd 9529: out = 12'h98F;
            14'd 9530: out = 12'h990;
            14'd 9531: out = 12'h990;
            14'd 9532: out = 12'h991;
            14'd 9533: out = 12'h991;
            14'd 9534: out = 12'h991;
            14'd 9535: out = 12'h992;
            14'd 9536: out = 12'h992;
            14'd 9537: out = 12'h992;
            14'd 9538: out = 12'h993;
            14'd 9539: out = 12'h993;
            14'd 9540: out = 12'h993;
            14'd 9541: out = 12'h994;
            14'd 9542: out = 12'h994;
            14'd 9543: out = 12'h994;
            14'd 9544: out = 12'h995;
            14'd 9545: out = 12'h995;
            14'd 9546: out = 12'h996;
            14'd 9547: out = 12'h996;
            14'd 9548: out = 12'h996;
            14'd 9549: out = 12'h997;
            14'd 9550: out = 12'h997;
            14'd 9551: out = 12'h997;
            14'd 9552: out = 12'h998;
            14'd 9553: out = 12'h998;
            14'd 9554: out = 12'h998;
            14'd 9555: out = 12'h999;
            14'd 9556: out = 12'h999;
            14'd 9557: out = 12'h999;
            14'd 9558: out = 12'h99A;
            14'd 9559: out = 12'h99A;
            14'd 9560: out = 12'h99B;
            14'd 9561: out = 12'h99B;
            14'd 9562: out = 12'h99B;
            14'd 9563: out = 12'h99C;
            14'd 9564: out = 12'h99C;
            14'd 9565: out = 12'h99C;
            14'd 9566: out = 12'h99D;
            14'd 9567: out = 12'h99D;
            14'd 9568: out = 12'h99D;
            14'd 9569: out = 12'h99E;
            14'd 9570: out = 12'h99E;
            14'd 9571: out = 12'h99F;
            14'd 9572: out = 12'h99F;
            14'd 9573: out = 12'h99F;
            14'd 9574: out = 12'h9A0;
            14'd 9575: out = 12'h9A0;
            14'd 9576: out = 12'h9A0;
            14'd 9577: out = 12'h9A1;
            14'd 9578: out = 12'h9A1;
            14'd 9579: out = 12'h9A1;
            14'd 9580: out = 12'h9A2;
            14'd 9581: out = 12'h9A2;
            14'd 9582: out = 12'h9A3;
            14'd 9583: out = 12'h9A3;
            14'd 9584: out = 12'h9A3;
            14'd 9585: out = 12'h9A4;
            14'd 9586: out = 12'h9A4;
            14'd 9587: out = 12'h9A4;
            14'd 9588: out = 12'h9A5;
            14'd 9589: out = 12'h9A5;
            14'd 9590: out = 12'h9A5;
            14'd 9591: out = 12'h9A6;
            14'd 9592: out = 12'h9A6;
            14'd 9593: out = 12'h9A7;
            14'd 9594: out = 12'h9A7;
            14'd 9595: out = 12'h9A7;
            14'd 9596: out = 12'h9A8;
            14'd 9597: out = 12'h9A8;
            14'd 9598: out = 12'h9A8;
            14'd 9599: out = 12'h9A9;
            14'd 9600: out = 12'h9A9;
            14'd 9601: out = 12'h9A9;
            14'd 9602: out = 12'h9AA;
            14'd 9603: out = 12'h9AA;
            14'd 9604: out = 12'h9AB;
            14'd 9605: out = 12'h9AB;
            14'd 9606: out = 12'h9AB;
            14'd 9607: out = 12'h9AC;
            14'd 9608: out = 12'h9AC;
            14'd 9609: out = 12'h9AC;
            14'd 9610: out = 12'h9AD;
            14'd 9611: out = 12'h9AD;
            14'd 9612: out = 12'h9AD;
            14'd 9613: out = 12'h9AE;
            14'd 9614: out = 12'h9AE;
            14'd 9615: out = 12'h9AF;
            14'd 9616: out = 12'h9AF;
            14'd 9617: out = 12'h9AF;
            14'd 9618: out = 12'h9B0;
            14'd 9619: out = 12'h9B0;
            14'd 9620: out = 12'h9B0;
            14'd 9621: out = 12'h9B1;
            14'd 9622: out = 12'h9B1;
            14'd 9623: out = 12'h9B1;
            14'd 9624: out = 12'h9B2;
            14'd 9625: out = 12'h9B2;
            14'd 9626: out = 12'h9B3;
            14'd 9627: out = 12'h9B3;
            14'd 9628: out = 12'h9B3;
            14'd 9629: out = 12'h9B4;
            14'd 9630: out = 12'h9B4;
            14'd 9631: out = 12'h9B4;
            14'd 9632: out = 12'h9B5;
            14'd 9633: out = 12'h9B5;
            14'd 9634: out = 12'h9B6;
            14'd 9635: out = 12'h9B6;
            14'd 9636: out = 12'h9B6;
            14'd 9637: out = 12'h9B7;
            14'd 9638: out = 12'h9B7;
            14'd 9639: out = 12'h9B7;
            14'd 9640: out = 12'h9B8;
            14'd 9641: out = 12'h9B8;
            14'd 9642: out = 12'h9B8;
            14'd 9643: out = 12'h9B9;
            14'd 9644: out = 12'h9B9;
            14'd 9645: out = 12'h9BA;
            14'd 9646: out = 12'h9BA;
            14'd 9647: out = 12'h9BA;
            14'd 9648: out = 12'h9BB;
            14'd 9649: out = 12'h9BB;
            14'd 9650: out = 12'h9BB;
            14'd 9651: out = 12'h9BC;
            14'd 9652: out = 12'h9BC;
            14'd 9653: out = 12'h9BD;
            14'd 9654: out = 12'h9BD;
            14'd 9655: out = 12'h9BD;
            14'd 9656: out = 12'h9BE;
            14'd 9657: out = 12'h9BE;
            14'd 9658: out = 12'h9BE;
            14'd 9659: out = 12'h9BF;
            14'd 9660: out = 12'h9BF;
            14'd 9661: out = 12'h9BF;
            14'd 9662: out = 12'h9C0;
            14'd 9663: out = 12'h9C0;
            14'd 9664: out = 12'h9C1;
            14'd 9665: out = 12'h9C1;
            14'd 9666: out = 12'h9C1;
            14'd 9667: out = 12'h9C2;
            14'd 9668: out = 12'h9C2;
            14'd 9669: out = 12'h9C2;
            14'd 9670: out = 12'h9C3;
            14'd 9671: out = 12'h9C3;
            14'd 9672: out = 12'h9C4;
            14'd 9673: out = 12'h9C4;
            14'd 9674: out = 12'h9C4;
            14'd 9675: out = 12'h9C5;
            14'd 9676: out = 12'h9C5;
            14'd 9677: out = 12'h9C5;
            14'd 9678: out = 12'h9C6;
            14'd 9679: out = 12'h9C6;
            14'd 9680: out = 12'h9C7;
            14'd 9681: out = 12'h9C7;
            14'd 9682: out = 12'h9C7;
            14'd 9683: out = 12'h9C8;
            14'd 9684: out = 12'h9C8;
            14'd 9685: out = 12'h9C8;
            14'd 9686: out = 12'h9C9;
            14'd 9687: out = 12'h9C9;
            14'd 9688: out = 12'h9CA;
            14'd 9689: out = 12'h9CA;
            14'd 9690: out = 12'h9CA;
            14'd 9691: out = 12'h9CB;
            14'd 9692: out = 12'h9CB;
            14'd 9693: out = 12'h9CB;
            14'd 9694: out = 12'h9CC;
            14'd 9695: out = 12'h9CC;
            14'd 9696: out = 12'h9CD;
            14'd 9697: out = 12'h9CD;
            14'd 9698: out = 12'h9CD;
            14'd 9699: out = 12'h9CE;
            14'd 9700: out = 12'h9CE;
            14'd 9701: out = 12'h9CE;
            14'd 9702: out = 12'h9CF;
            14'd 9703: out = 12'h9CF;
            14'd 9704: out = 12'h9D0;
            14'd 9705: out = 12'h9D0;
            14'd 9706: out = 12'h9D0;
            14'd 9707: out = 12'h9D1;
            14'd 9708: out = 12'h9D1;
            14'd 9709: out = 12'h9D1;
            14'd 9710: out = 12'h9D2;
            14'd 9711: out = 12'h9D2;
            14'd 9712: out = 12'h9D3;
            14'd 9713: out = 12'h9D3;
            14'd 9714: out = 12'h9D3;
            14'd 9715: out = 12'h9D4;
            14'd 9716: out = 12'h9D4;
            14'd 9717: out = 12'h9D4;
            14'd 9718: out = 12'h9D5;
            14'd 9719: out = 12'h9D5;
            14'd 9720: out = 12'h9D6;
            14'd 9721: out = 12'h9D6;
            14'd 9722: out = 12'h9D6;
            14'd 9723: out = 12'h9D7;
            14'd 9724: out = 12'h9D7;
            14'd 9725: out = 12'h9D7;
            14'd 9726: out = 12'h9D8;
            14'd 9727: out = 12'h9D8;
            14'd 9728: out = 12'h9D9;
            14'd 9729: out = 12'h9D9;
            14'd 9730: out = 12'h9D9;
            14'd 9731: out = 12'h9DA;
            14'd 9732: out = 12'h9DA;
            14'd 9733: out = 12'h9DB;
            14'd 9734: out = 12'h9DB;
            14'd 9735: out = 12'h9DB;
            14'd 9736: out = 12'h9DC;
            14'd 9737: out = 12'h9DC;
            14'd 9738: out = 12'h9DC;
            14'd 9739: out = 12'h9DD;
            14'd 9740: out = 12'h9DD;
            14'd 9741: out = 12'h9DE;
            14'd 9742: out = 12'h9DE;
            14'd 9743: out = 12'h9DE;
            14'd 9744: out = 12'h9DF;
            14'd 9745: out = 12'h9DF;
            14'd 9746: out = 12'h9DF;
            14'd 9747: out = 12'h9E0;
            14'd 9748: out = 12'h9E0;
            14'd 9749: out = 12'h9E1;
            14'd 9750: out = 12'h9E1;
            14'd 9751: out = 12'h9E1;
            14'd 9752: out = 12'h9E2;
            14'd 9753: out = 12'h9E2;
            14'd 9754: out = 12'h9E3;
            14'd 9755: out = 12'h9E3;
            14'd 9756: out = 12'h9E3;
            14'd 9757: out = 12'h9E4;
            14'd 9758: out = 12'h9E4;
            14'd 9759: out = 12'h9E4;
            14'd 9760: out = 12'h9E5;
            14'd 9761: out = 12'h9E5;
            14'd 9762: out = 12'h9E6;
            14'd 9763: out = 12'h9E6;
            14'd 9764: out = 12'h9E6;
            14'd 9765: out = 12'h9E7;
            14'd 9766: out = 12'h9E7;
            14'd 9767: out = 12'h9E7;
            14'd 9768: out = 12'h9E8;
            14'd 9769: out = 12'h9E8;
            14'd 9770: out = 12'h9E9;
            14'd 9771: out = 12'h9E9;
            14'd 9772: out = 12'h9E9;
            14'd 9773: out = 12'h9EA;
            14'd 9774: out = 12'h9EA;
            14'd 9775: out = 12'h9EB;
            14'd 9776: out = 12'h9EB;
            14'd 9777: out = 12'h9EB;
            14'd 9778: out = 12'h9EC;
            14'd 9779: out = 12'h9EC;
            14'd 9780: out = 12'h9EC;
            14'd 9781: out = 12'h9ED;
            14'd 9782: out = 12'h9ED;
            14'd 9783: out = 12'h9EE;
            14'd 9784: out = 12'h9EE;
            14'd 9785: out = 12'h9EE;
            14'd 9786: out = 12'h9EF;
            14'd 9787: out = 12'h9EF;
            14'd 9788: out = 12'h9F0;
            14'd 9789: out = 12'h9F0;
            14'd 9790: out = 12'h9F0;
            14'd 9791: out = 12'h9F1;
            14'd 9792: out = 12'h9F1;
            14'd 9793: out = 12'h9F1;
            14'd 9794: out = 12'h9F2;
            14'd 9795: out = 12'h9F2;
            14'd 9796: out = 12'h9F3;
            14'd 9797: out = 12'h9F3;
            14'd 9798: out = 12'h9F3;
            14'd 9799: out = 12'h9F4;
            14'd 9800: out = 12'h9F4;
            14'd 9801: out = 12'h9F5;
            14'd 9802: out = 12'h9F5;
            14'd 9803: out = 12'h9F5;
            14'd 9804: out = 12'h9F6;
            14'd 9805: out = 12'h9F6;
            14'd 9806: out = 12'h9F7;
            14'd 9807: out = 12'h9F7;
            14'd 9808: out = 12'h9F7;
            14'd 9809: out = 12'h9F8;
            14'd 9810: out = 12'h9F8;
            14'd 9811: out = 12'h9F8;
            14'd 9812: out = 12'h9F9;
            14'd 9813: out = 12'h9F9;
            14'd 9814: out = 12'h9FA;
            14'd 9815: out = 12'h9FA;
            14'd 9816: out = 12'h9FA;
            14'd 9817: out = 12'h9FB;
            14'd 9818: out = 12'h9FB;
            14'd 9819: out = 12'h9FC;
            14'd 9820: out = 12'h9FC;
            14'd 9821: out = 12'h9FC;
            14'd 9822: out = 12'h9FD;
            14'd 9823: out = 12'h9FD;
            14'd 9824: out = 12'h9FE;
            14'd 9825: out = 12'h9FE;
            14'd 9826: out = 12'h9FE;
            14'd 9827: out = 12'h9FF;
            14'd 9828: out = 12'h9FF;
            14'd 9829: out = 12'h9FF;
            14'd 9830: out = 12'hA00;
            14'd 9831: out = 12'hA00;
            14'd 9832: out = 12'hA01;
            14'd 9833: out = 12'hA01;
            14'd 9834: out = 12'hA01;
            14'd 9835: out = 12'hA02;
            14'd 9836: out = 12'hA02;
            14'd 9837: out = 12'hA03;
            14'd 9838: out = 12'hA03;
            14'd 9839: out = 12'hA03;
            14'd 9840: out = 12'hA04;
            14'd 9841: out = 12'hA04;
            14'd 9842: out = 12'hA05;
            14'd 9843: out = 12'hA05;
            14'd 9844: out = 12'hA05;
            14'd 9845: out = 12'hA06;
            14'd 9846: out = 12'hA06;
            14'd 9847: out = 12'hA07;
            14'd 9848: out = 12'hA07;
            14'd 9849: out = 12'hA07;
            14'd 9850: out = 12'hA08;
            14'd 9851: out = 12'hA08;
            14'd 9852: out = 12'hA08;
            14'd 9853: out = 12'hA09;
            14'd 9854: out = 12'hA09;
            14'd 9855: out = 12'hA0A;
            14'd 9856: out = 12'hA0A;
            14'd 9857: out = 12'hA0A;
            14'd 9858: out = 12'hA0B;
            14'd 9859: out = 12'hA0B;
            14'd 9860: out = 12'hA0C;
            14'd 9861: out = 12'hA0C;
            14'd 9862: out = 12'hA0C;
            14'd 9863: out = 12'hA0D;
            14'd 9864: out = 12'hA0D;
            14'd 9865: out = 12'hA0E;
            14'd 9866: out = 12'hA0E;
            14'd 9867: out = 12'hA0E;
            14'd 9868: out = 12'hA0F;
            14'd 9869: out = 12'hA0F;
            14'd 9870: out = 12'hA10;
            14'd 9871: out = 12'hA10;
            14'd 9872: out = 12'hA10;
            14'd 9873: out = 12'hA11;
            14'd 9874: out = 12'hA11;
            14'd 9875: out = 12'hA12;
            14'd 9876: out = 12'hA12;
            14'd 9877: out = 12'hA12;
            14'd 9878: out = 12'hA13;
            14'd 9879: out = 12'hA13;
            14'd 9880: out = 12'hA14;
            14'd 9881: out = 12'hA14;
            14'd 9882: out = 12'hA14;
            14'd 9883: out = 12'hA15;
            14'd 9884: out = 12'hA15;
            14'd 9885: out = 12'hA16;
            14'd 9886: out = 12'hA16;
            14'd 9887: out = 12'hA16;
            14'd 9888: out = 12'hA17;
            14'd 9889: out = 12'hA17;
            14'd 9890: out = 12'hA17;
            14'd 9891: out = 12'hA18;
            14'd 9892: out = 12'hA18;
            14'd 9893: out = 12'hA19;
            14'd 9894: out = 12'hA19;
            14'd 9895: out = 12'hA19;
            14'd 9896: out = 12'hA1A;
            14'd 9897: out = 12'hA1A;
            14'd 9898: out = 12'hA1B;
            14'd 9899: out = 12'hA1B;
            14'd 9900: out = 12'hA1B;
            14'd 9901: out = 12'hA1C;
            14'd 9902: out = 12'hA1C;
            14'd 9903: out = 12'hA1D;
            14'd 9904: out = 12'hA1D;
            14'd 9905: out = 12'hA1D;
            14'd 9906: out = 12'hA1E;
            14'd 9907: out = 12'hA1E;
            14'd 9908: out = 12'hA1F;
            14'd 9909: out = 12'hA1F;
            14'd 9910: out = 12'hA1F;
            14'd 9911: out = 12'hA20;
            14'd 9912: out = 12'hA20;
            14'd 9913: out = 12'hA21;
            14'd 9914: out = 12'hA21;
            14'd 9915: out = 12'hA21;
            14'd 9916: out = 12'hA22;
            14'd 9917: out = 12'hA22;
            14'd 9918: out = 12'hA23;
            14'd 9919: out = 12'hA23;
            14'd 9920: out = 12'hA23;
            14'd 9921: out = 12'hA24;
            14'd 9922: out = 12'hA24;
            14'd 9923: out = 12'hA25;
            14'd 9924: out = 12'hA25;
            14'd 9925: out = 12'hA25;
            14'd 9926: out = 12'hA26;
            14'd 9927: out = 12'hA26;
            14'd 9928: out = 12'hA27;
            14'd 9929: out = 12'hA27;
            14'd 9930: out = 12'hA28;
            14'd 9931: out = 12'hA28;
            14'd 9932: out = 12'hA28;
            14'd 9933: out = 12'hA29;
            14'd 9934: out = 12'hA29;
            14'd 9935: out = 12'hA2A;
            14'd 9936: out = 12'hA2A;
            14'd 9937: out = 12'hA2A;
            14'd 9938: out = 12'hA2B;
            14'd 9939: out = 12'hA2B;
            14'd 9940: out = 12'hA2C;
            14'd 9941: out = 12'hA2C;
            14'd 9942: out = 12'hA2C;
            14'd 9943: out = 12'hA2D;
            14'd 9944: out = 12'hA2D;
            14'd 9945: out = 12'hA2E;
            14'd 9946: out = 12'hA2E;
            14'd 9947: out = 12'hA2E;
            14'd 9948: out = 12'hA2F;
            14'd 9949: out = 12'hA2F;
            14'd 9950: out = 12'hA30;
            14'd 9951: out = 12'hA30;
            14'd 9952: out = 12'hA30;
            14'd 9953: out = 12'hA31;
            14'd 9954: out = 12'hA31;
            14'd 9955: out = 12'hA32;
            14'd 9956: out = 12'hA32;
            14'd 9957: out = 12'hA32;
            14'd 9958: out = 12'hA33;
            14'd 9959: out = 12'hA33;
            14'd 9960: out = 12'hA34;
            14'd 9961: out = 12'hA34;
            14'd 9962: out = 12'hA34;
            14'd 9963: out = 12'hA35;
            14'd 9964: out = 12'hA35;
            14'd 9965: out = 12'hA36;
            14'd 9966: out = 12'hA36;
            14'd 9967: out = 12'hA36;
            14'd 9968: out = 12'hA37;
            14'd 9969: out = 12'hA37;
            14'd 9970: out = 12'hA38;
            14'd 9971: out = 12'hA38;
            14'd 9972: out = 12'hA39;
            14'd 9973: out = 12'hA39;
            14'd 9974: out = 12'hA39;
            14'd 9975: out = 12'hA3A;
            14'd 9976: out = 12'hA3A;
            14'd 9977: out = 12'hA3B;
            14'd 9978: out = 12'hA3B;
            14'd 9979: out = 12'hA3B;
            14'd 9980: out = 12'hA3C;
            14'd 9981: out = 12'hA3C;
            14'd 9982: out = 12'hA3D;
            14'd 9983: out = 12'hA3D;
            14'd 9984: out = 12'hA3D;
            14'd 9985: out = 12'hA3E;
            14'd 9986: out = 12'hA3E;
            14'd 9987: out = 12'hA3F;
            14'd 9988: out = 12'hA3F;
            14'd 9989: out = 12'hA3F;
            14'd 9990: out = 12'hA40;
            14'd 9991: out = 12'hA40;
            14'd 9992: out = 12'hA41;
            14'd 9993: out = 12'hA41;
            14'd 9994: out = 12'hA42;
            14'd 9995: out = 12'hA42;
            14'd 9996: out = 12'hA42;
            14'd 9997: out = 12'hA43;
            14'd 9998: out = 12'hA43;
            14'd 9999: out = 12'hA44;
            14'd10000: out = 12'hA44;
            14'd10001: out = 12'hA44;
            14'd10002: out = 12'hA45;
            14'd10003: out = 12'hA45;
            14'd10004: out = 12'hA46;
            14'd10005: out = 12'hA46;
            14'd10006: out = 12'hA46;
            14'd10007: out = 12'hA47;
            14'd10008: out = 12'hA47;
            14'd10009: out = 12'hA48;
            14'd10010: out = 12'hA48;
            14'd10011: out = 12'hA49;
            14'd10012: out = 12'hA49;
            14'd10013: out = 12'hA49;
            14'd10014: out = 12'hA4A;
            14'd10015: out = 12'hA4A;
            14'd10016: out = 12'hA4B;
            14'd10017: out = 12'hA4B;
            14'd10018: out = 12'hA4B;
            14'd10019: out = 12'hA4C;
            14'd10020: out = 12'hA4C;
            14'd10021: out = 12'hA4D;
            14'd10022: out = 12'hA4D;
            14'd10023: out = 12'hA4E;
            14'd10024: out = 12'hA4E;
            14'd10025: out = 12'hA4E;
            14'd10026: out = 12'hA4F;
            14'd10027: out = 12'hA4F;
            14'd10028: out = 12'hA50;
            14'd10029: out = 12'hA50;
            14'd10030: out = 12'hA50;
            14'd10031: out = 12'hA51;
            14'd10032: out = 12'hA51;
            14'd10033: out = 12'hA52;
            14'd10034: out = 12'hA52;
            14'd10035: out = 12'hA52;
            14'd10036: out = 12'hA53;
            14'd10037: out = 12'hA53;
            14'd10038: out = 12'hA54;
            14'd10039: out = 12'hA54;
            14'd10040: out = 12'hA55;
            14'd10041: out = 12'hA55;
            14'd10042: out = 12'hA55;
            14'd10043: out = 12'hA56;
            14'd10044: out = 12'hA56;
            14'd10045: out = 12'hA57;
            14'd10046: out = 12'hA57;
            14'd10047: out = 12'hA58;
            14'd10048: out = 12'hA58;
            14'd10049: out = 12'hA58;
            14'd10050: out = 12'hA59;
            14'd10051: out = 12'hA59;
            14'd10052: out = 12'hA5A;
            14'd10053: out = 12'hA5A;
            14'd10054: out = 12'hA5A;
            14'd10055: out = 12'hA5B;
            14'd10056: out = 12'hA5B;
            14'd10057: out = 12'hA5C;
            14'd10058: out = 12'hA5C;
            14'd10059: out = 12'hA5D;
            14'd10060: out = 12'hA5D;
            14'd10061: out = 12'hA5D;
            14'd10062: out = 12'hA5E;
            14'd10063: out = 12'hA5E;
            14'd10064: out = 12'hA5F;
            14'd10065: out = 12'hA5F;
            14'd10066: out = 12'hA5F;
            14'd10067: out = 12'hA60;
            14'd10068: out = 12'hA60;
            14'd10069: out = 12'hA61;
            14'd10070: out = 12'hA61;
            14'd10071: out = 12'hA62;
            14'd10072: out = 12'hA62;
            14'd10073: out = 12'hA62;
            14'd10074: out = 12'hA63;
            14'd10075: out = 12'hA63;
            14'd10076: out = 12'hA64;
            14'd10077: out = 12'hA64;
            14'd10078: out = 12'hA65;
            14'd10079: out = 12'hA65;
            14'd10080: out = 12'hA65;
            14'd10081: out = 12'hA66;
            14'd10082: out = 12'hA66;
            14'd10083: out = 12'hA67;
            14'd10084: out = 12'hA67;
            14'd10085: out = 12'hA67;
            14'd10086: out = 12'hA68;
            14'd10087: out = 12'hA68;
            14'd10088: out = 12'hA69;
            14'd10089: out = 12'hA69;
            14'd10090: out = 12'hA6A;
            14'd10091: out = 12'hA6A;
            14'd10092: out = 12'hA6A;
            14'd10093: out = 12'hA6B;
            14'd10094: out = 12'hA6B;
            14'd10095: out = 12'hA6C;
            14'd10096: out = 12'hA6C;
            14'd10097: out = 12'hA6D;
            14'd10098: out = 12'hA6D;
            14'd10099: out = 12'hA6D;
            14'd10100: out = 12'hA6E;
            14'd10101: out = 12'hA6E;
            14'd10102: out = 12'hA6F;
            14'd10103: out = 12'hA6F;
            14'd10104: out = 12'hA70;
            14'd10105: out = 12'hA70;
            14'd10106: out = 12'hA70;
            14'd10107: out = 12'hA71;
            14'd10108: out = 12'hA71;
            14'd10109: out = 12'hA72;
            14'd10110: out = 12'hA72;
            14'd10111: out = 12'hA73;
            14'd10112: out = 12'hA73;
            14'd10113: out = 12'hA73;
            14'd10114: out = 12'hA74;
            14'd10115: out = 12'hA74;
            14'd10116: out = 12'hA75;
            14'd10117: out = 12'hA75;
            14'd10118: out = 12'hA76;
            14'd10119: out = 12'hA76;
            14'd10120: out = 12'hA76;
            14'd10121: out = 12'hA77;
            14'd10122: out = 12'hA77;
            14'd10123: out = 12'hA78;
            14'd10124: out = 12'hA78;
            14'd10125: out = 12'hA78;
            14'd10126: out = 12'hA79;
            14'd10127: out = 12'hA79;
            14'd10128: out = 12'hA7A;
            14'd10129: out = 12'hA7A;
            14'd10130: out = 12'hA7B;
            14'd10131: out = 12'hA7B;
            14'd10132: out = 12'hA7B;
            14'd10133: out = 12'hA7C;
            14'd10134: out = 12'hA7C;
            14'd10135: out = 12'hA7D;
            14'd10136: out = 12'hA7D;
            14'd10137: out = 12'hA7E;
            14'd10138: out = 12'hA7E;
            14'd10139: out = 12'hA7F;
            14'd10140: out = 12'hA7F;
            14'd10141: out = 12'hA7F;
            14'd10142: out = 12'hA80;
            14'd10143: out = 12'hA80;
            14'd10144: out = 12'hA81;
            14'd10145: out = 12'hA81;
            14'd10146: out = 12'hA82;
            14'd10147: out = 12'hA82;
            14'd10148: out = 12'hA82;
            14'd10149: out = 12'hA83;
            14'd10150: out = 12'hA83;
            14'd10151: out = 12'hA84;
            14'd10152: out = 12'hA84;
            14'd10153: out = 12'hA85;
            14'd10154: out = 12'hA85;
            14'd10155: out = 12'hA85;
            14'd10156: out = 12'hA86;
            14'd10157: out = 12'hA86;
            14'd10158: out = 12'hA87;
            14'd10159: out = 12'hA87;
            14'd10160: out = 12'hA88;
            14'd10161: out = 12'hA88;
            14'd10162: out = 12'hA88;
            14'd10163: out = 12'hA89;
            14'd10164: out = 12'hA89;
            14'd10165: out = 12'hA8A;
            14'd10166: out = 12'hA8A;
            14'd10167: out = 12'hA8B;
            14'd10168: out = 12'hA8B;
            14'd10169: out = 12'hA8B;
            14'd10170: out = 12'hA8C;
            14'd10171: out = 12'hA8C;
            14'd10172: out = 12'hA8D;
            14'd10173: out = 12'hA8D;
            14'd10174: out = 12'hA8E;
            14'd10175: out = 12'hA8E;
            14'd10176: out = 12'hA8F;
            14'd10177: out = 12'hA8F;
            14'd10178: out = 12'hA8F;
            14'd10179: out = 12'hA90;
            14'd10180: out = 12'hA90;
            14'd10181: out = 12'hA91;
            14'd10182: out = 12'hA91;
            14'd10183: out = 12'hA92;
            14'd10184: out = 12'hA92;
            14'd10185: out = 12'hA92;
            14'd10186: out = 12'hA93;
            14'd10187: out = 12'hA93;
            14'd10188: out = 12'hA94;
            14'd10189: out = 12'hA94;
            14'd10190: out = 12'hA95;
            14'd10191: out = 12'hA95;
            14'd10192: out = 12'hA95;
            14'd10193: out = 12'hA96;
            14'd10194: out = 12'hA96;
            14'd10195: out = 12'hA97;
            14'd10196: out = 12'hA97;
            14'd10197: out = 12'hA98;
            14'd10198: out = 12'hA98;
            14'd10199: out = 12'hA99;
            14'd10200: out = 12'hA99;
            14'd10201: out = 12'hA99;
            14'd10202: out = 12'hA9A;
            14'd10203: out = 12'hA9A;
            14'd10204: out = 12'hA9B;
            14'd10205: out = 12'hA9B;
            14'd10206: out = 12'hA9C;
            14'd10207: out = 12'hA9C;
            14'd10208: out = 12'hA9D;
            14'd10209: out = 12'hA9D;
            14'd10210: out = 12'hA9D;
            14'd10211: out = 12'hA9E;
            14'd10212: out = 12'hA9E;
            14'd10213: out = 12'hA9F;
            14'd10214: out = 12'hA9F;
            14'd10215: out = 12'hAA0;
            14'd10216: out = 12'hAA0;
            14'd10217: out = 12'hAA0;
            14'd10218: out = 12'hAA1;
            14'd10219: out = 12'hAA1;
            14'd10220: out = 12'hAA2;
            14'd10221: out = 12'hAA2;
            14'd10222: out = 12'hAA3;
            14'd10223: out = 12'hAA3;
            14'd10224: out = 12'hAA4;
            14'd10225: out = 12'hAA4;
            14'd10226: out = 12'hAA4;
            14'd10227: out = 12'hAA5;
            14'd10228: out = 12'hAA5;
            14'd10229: out = 12'hAA6;
            14'd10230: out = 12'hAA6;
            14'd10231: out = 12'hAA7;
            14'd10232: out = 12'hAA7;
            14'd10233: out = 12'hAA8;
            14'd10234: out = 12'hAA8;
            14'd10235: out = 12'hAA8;
            14'd10236: out = 12'hAA9;
            14'd10237: out = 12'hAA9;
            14'd10238: out = 12'hAAA;
            14'd10239: out = 12'hAAA;
            14'd10240: out = 12'hAAB;
            14'd10241: out = 12'hAAB;
            14'd10242: out = 12'hAAC;
            14'd10243: out = 12'hAAC;
            14'd10244: out = 12'hAAC;
            14'd10245: out = 12'hAAD;
            14'd10246: out = 12'hAAD;
            14'd10247: out = 12'hAAE;
            14'd10248: out = 12'hAAE;
            14'd10249: out = 12'hAAF;
            14'd10250: out = 12'hAAF;
            14'd10251: out = 12'hAB0;
            14'd10252: out = 12'hAB0;
            14'd10253: out = 12'hAB0;
            14'd10254: out = 12'hAB1;
            14'd10255: out = 12'hAB1;
            14'd10256: out = 12'hAB2;
            14'd10257: out = 12'hAB2;
            14'd10258: out = 12'hAB3;
            14'd10259: out = 12'hAB3;
            14'd10260: out = 12'hAB4;
            14'd10261: out = 12'hAB4;
            14'd10262: out = 12'hAB4;
            14'd10263: out = 12'hAB5;
            14'd10264: out = 12'hAB5;
            14'd10265: out = 12'hAB6;
            14'd10266: out = 12'hAB6;
            14'd10267: out = 12'hAB7;
            14'd10268: out = 12'hAB7;
            14'd10269: out = 12'hAB8;
            14'd10270: out = 12'hAB8;
            14'd10271: out = 12'hAB9;
            14'd10272: out = 12'hAB9;
            14'd10273: out = 12'hAB9;
            14'd10274: out = 12'hABA;
            14'd10275: out = 12'hABA;
            14'd10276: out = 12'hABB;
            14'd10277: out = 12'hABB;
            14'd10278: out = 12'hABC;
            14'd10279: out = 12'hABC;
            14'd10280: out = 12'hABD;
            14'd10281: out = 12'hABD;
            14'd10282: out = 12'hABD;
            14'd10283: out = 12'hABE;
            14'd10284: out = 12'hABE;
            14'd10285: out = 12'hABF;
            14'd10286: out = 12'hABF;
            14'd10287: out = 12'hAC0;
            14'd10288: out = 12'hAC0;
            14'd10289: out = 12'hAC1;
            14'd10290: out = 12'hAC1;
            14'd10291: out = 12'hAC2;
            14'd10292: out = 12'hAC2;
            14'd10293: out = 12'hAC2;
            14'd10294: out = 12'hAC3;
            14'd10295: out = 12'hAC3;
            14'd10296: out = 12'hAC4;
            14'd10297: out = 12'hAC4;
            14'd10298: out = 12'hAC5;
            14'd10299: out = 12'hAC5;
            14'd10300: out = 12'hAC6;
            14'd10301: out = 12'hAC6;
            14'd10302: out = 12'hAC7;
            14'd10303: out = 12'hAC7;
            14'd10304: out = 12'hAC7;
            14'd10305: out = 12'hAC8;
            14'd10306: out = 12'hAC8;
            14'd10307: out = 12'hAC9;
            14'd10308: out = 12'hAC9;
            14'd10309: out = 12'hACA;
            14'd10310: out = 12'hACA;
            14'd10311: out = 12'hACB;
            14'd10312: out = 12'hACB;
            14'd10313: out = 12'hACC;
            14'd10314: out = 12'hACC;
            14'd10315: out = 12'hACC;
            14'd10316: out = 12'hACD;
            14'd10317: out = 12'hACD;
            14'd10318: out = 12'hACE;
            14'd10319: out = 12'hACE;
            14'd10320: out = 12'hACF;
            14'd10321: out = 12'hACF;
            14'd10322: out = 12'hAD0;
            14'd10323: out = 12'hAD0;
            14'd10324: out = 12'hAD1;
            14'd10325: out = 12'hAD1;
            14'd10326: out = 12'hAD1;
            14'd10327: out = 12'hAD2;
            14'd10328: out = 12'hAD2;
            14'd10329: out = 12'hAD3;
            14'd10330: out = 12'hAD3;
            14'd10331: out = 12'hAD4;
            14'd10332: out = 12'hAD4;
            14'd10333: out = 12'hAD5;
            14'd10334: out = 12'hAD5;
            14'd10335: out = 12'hAD6;
            14'd10336: out = 12'hAD6;
            14'd10337: out = 12'hAD6;
            14'd10338: out = 12'hAD7;
            14'd10339: out = 12'hAD7;
            14'd10340: out = 12'hAD8;
            14'd10341: out = 12'hAD8;
            14'd10342: out = 12'hAD9;
            14'd10343: out = 12'hAD9;
            14'd10344: out = 12'hADA;
            14'd10345: out = 12'hADA;
            14'd10346: out = 12'hADB;
            14'd10347: out = 12'hADB;
            14'd10348: out = 12'hADC;
            14'd10349: out = 12'hADC;
            14'd10350: out = 12'hADC;
            14'd10351: out = 12'hADD;
            14'd10352: out = 12'hADD;
            14'd10353: out = 12'hADE;
            14'd10354: out = 12'hADE;
            14'd10355: out = 12'hADF;
            14'd10356: out = 12'hADF;
            14'd10357: out = 12'hAE0;
            14'd10358: out = 12'hAE0;
            14'd10359: out = 12'hAE1;
            14'd10360: out = 12'hAE1;
            14'd10361: out = 12'hAE2;
            14'd10362: out = 12'hAE2;
            14'd10363: out = 12'hAE2;
            14'd10364: out = 12'hAE3;
            14'd10365: out = 12'hAE3;
            14'd10366: out = 12'hAE4;
            14'd10367: out = 12'hAE4;
            14'd10368: out = 12'hAE5;
            14'd10369: out = 12'hAE5;
            14'd10370: out = 12'hAE6;
            14'd10371: out = 12'hAE6;
            14'd10372: out = 12'hAE7;
            14'd10373: out = 12'hAE7;
            14'd10374: out = 12'hAE8;
            14'd10375: out = 12'hAE8;
            14'd10376: out = 12'hAE8;
            14'd10377: out = 12'hAE9;
            14'd10378: out = 12'hAE9;
            14'd10379: out = 12'hAEA;
            14'd10380: out = 12'hAEA;
            14'd10381: out = 12'hAEB;
            14'd10382: out = 12'hAEB;
            14'd10383: out = 12'hAEC;
            14'd10384: out = 12'hAEC;
            14'd10385: out = 12'hAED;
            14'd10386: out = 12'hAED;
            14'd10387: out = 12'hAEE;
            14'd10388: out = 12'hAEE;
            14'd10389: out = 12'hAEF;
            14'd10390: out = 12'hAEF;
            14'd10391: out = 12'hAEF;
            14'd10392: out = 12'hAF0;
            14'd10393: out = 12'hAF0;
            14'd10394: out = 12'hAF1;
            14'd10395: out = 12'hAF1;
            14'd10396: out = 12'hAF2;
            14'd10397: out = 12'hAF2;
            14'd10398: out = 12'hAF3;
            14'd10399: out = 12'hAF3;
            14'd10400: out = 12'hAF4;
            14'd10401: out = 12'hAF4;
            14'd10402: out = 12'hAF5;
            14'd10403: out = 12'hAF5;
            14'd10404: out = 12'hAF6;
            14'd10405: out = 12'hAF6;
            14'd10406: out = 12'hAF6;
            14'd10407: out = 12'hAF7;
            14'd10408: out = 12'hAF7;
            14'd10409: out = 12'hAF8;
            14'd10410: out = 12'hAF8;
            14'd10411: out = 12'hAF9;
            14'd10412: out = 12'hAF9;
            14'd10413: out = 12'hAFA;
            14'd10414: out = 12'hAFA;
            14'd10415: out = 12'hAFB;
            14'd10416: out = 12'hAFB;
            14'd10417: out = 12'hAFC;
            14'd10418: out = 12'hAFC;
            14'd10419: out = 12'hAFD;
            14'd10420: out = 12'hAFD;
            14'd10421: out = 12'hAFE;
            14'd10422: out = 12'hAFE;
            14'd10423: out = 12'hAFE;
            14'd10424: out = 12'hAFF;
            14'd10425: out = 12'hAFF;
            14'd10426: out = 12'hB00;
            14'd10427: out = 12'hB00;
            14'd10428: out = 12'hB01;
            14'd10429: out = 12'hB01;
            14'd10430: out = 12'hB02;
            14'd10431: out = 12'hB02;
            14'd10432: out = 12'hB03;
            14'd10433: out = 12'hB03;
            14'd10434: out = 12'hB04;
            14'd10435: out = 12'hB04;
            14'd10436: out = 12'hB05;
            14'd10437: out = 12'hB05;
            14'd10438: out = 12'hB06;
            14'd10439: out = 12'hB06;
            14'd10440: out = 12'hB07;
            14'd10441: out = 12'hB07;
            14'd10442: out = 12'hB07;
            14'd10443: out = 12'hB08;
            14'd10444: out = 12'hB08;
            14'd10445: out = 12'hB09;
            14'd10446: out = 12'hB09;
            14'd10447: out = 12'hB0A;
            14'd10448: out = 12'hB0A;
            14'd10449: out = 12'hB0B;
            14'd10450: out = 12'hB0B;
            14'd10451: out = 12'hB0C;
            14'd10452: out = 12'hB0C;
            14'd10453: out = 12'hB0D;
            14'd10454: out = 12'hB0D;
            14'd10455: out = 12'hB0E;
            14'd10456: out = 12'hB0E;
            14'd10457: out = 12'hB0F;
            14'd10458: out = 12'hB0F;
            14'd10459: out = 12'hB10;
            14'd10460: out = 12'hB10;
            14'd10461: out = 12'hB11;
            14'd10462: out = 12'hB11;
            14'd10463: out = 12'hB12;
            14'd10464: out = 12'hB12;
            14'd10465: out = 12'hB12;
            14'd10466: out = 12'hB13;
            14'd10467: out = 12'hB13;
            14'd10468: out = 12'hB14;
            14'd10469: out = 12'hB14;
            14'd10470: out = 12'hB15;
            14'd10471: out = 12'hB15;
            14'd10472: out = 12'hB16;
            14'd10473: out = 12'hB16;
            14'd10474: out = 12'hB17;
            14'd10475: out = 12'hB17;
            14'd10476: out = 12'hB18;
            14'd10477: out = 12'hB18;
            14'd10478: out = 12'hB19;
            14'd10479: out = 12'hB19;
            14'd10480: out = 12'hB1A;
            14'd10481: out = 12'hB1A;
            14'd10482: out = 12'hB1B;
            14'd10483: out = 12'hB1B;
            14'd10484: out = 12'hB1C;
            14'd10485: out = 12'hB1C;
            14'd10486: out = 12'hB1D;
            14'd10487: out = 12'hB1D;
            14'd10488: out = 12'hB1E;
            14'd10489: out = 12'hB1E;
            14'd10490: out = 12'hB1E;
            14'd10491: out = 12'hB1F;
            14'd10492: out = 12'hB1F;
            14'd10493: out = 12'hB20;
            14'd10494: out = 12'hB20;
            14'd10495: out = 12'hB21;
            14'd10496: out = 12'hB21;
            14'd10497: out = 12'hB22;
            14'd10498: out = 12'hB22;
            14'd10499: out = 12'hB23;
            14'd10500: out = 12'hB23;
            14'd10501: out = 12'hB24;
            14'd10502: out = 12'hB24;
            14'd10503: out = 12'hB25;
            14'd10504: out = 12'hB25;
            14'd10505: out = 12'hB26;
            14'd10506: out = 12'hB26;
            14'd10507: out = 12'hB27;
            14'd10508: out = 12'hB27;
            14'd10509: out = 12'hB28;
            14'd10510: out = 12'hB28;
            14'd10511: out = 12'hB29;
            14'd10512: out = 12'hB29;
            14'd10513: out = 12'hB2A;
            14'd10514: out = 12'hB2A;
            14'd10515: out = 12'hB2B;
            14'd10516: out = 12'hB2B;
            14'd10517: out = 12'hB2C;
            14'd10518: out = 12'hB2C;
            14'd10519: out = 12'hB2D;
            14'd10520: out = 12'hB2D;
            14'd10521: out = 12'hB2E;
            14'd10522: out = 12'hB2E;
            14'd10523: out = 12'hB2F;
            14'd10524: out = 12'hB2F;
            14'd10525: out = 12'hB2F;
            14'd10526: out = 12'hB30;
            14'd10527: out = 12'hB30;
            14'd10528: out = 12'hB31;
            14'd10529: out = 12'hB31;
            14'd10530: out = 12'hB32;
            14'd10531: out = 12'hB32;
            14'd10532: out = 12'hB33;
            14'd10533: out = 12'hB33;
            14'd10534: out = 12'hB34;
            14'd10535: out = 12'hB34;
            14'd10536: out = 12'hB35;
            14'd10537: out = 12'hB35;
            14'd10538: out = 12'hB36;
            14'd10539: out = 12'hB36;
            14'd10540: out = 12'hB37;
            14'd10541: out = 12'hB37;
            14'd10542: out = 12'hB38;
            14'd10543: out = 12'hB38;
            14'd10544: out = 12'hB39;
            14'd10545: out = 12'hB39;
            14'd10546: out = 12'hB3A;
            14'd10547: out = 12'hB3A;
            14'd10548: out = 12'hB3B;
            14'd10549: out = 12'hB3B;
            14'd10550: out = 12'hB3C;
            14'd10551: out = 12'hB3C;
            14'd10552: out = 12'hB3D;
            14'd10553: out = 12'hB3D;
            14'd10554: out = 12'hB3E;
            14'd10555: out = 12'hB3E;
            14'd10556: out = 12'hB3F;
            14'd10557: out = 12'hB3F;
            14'd10558: out = 12'hB40;
            14'd10559: out = 12'hB40;
            14'd10560: out = 12'hB41;
            14'd10561: out = 12'hB41;
            14'd10562: out = 12'hB42;
            14'd10563: out = 12'hB42;
            14'd10564: out = 12'hB43;
            14'd10565: out = 12'hB43;
            14'd10566: out = 12'hB44;
            14'd10567: out = 12'hB44;
            14'd10568: out = 12'hB45;
            14'd10569: out = 12'hB45;
            14'd10570: out = 12'hB46;
            14'd10571: out = 12'hB46;
            14'd10572: out = 12'hB47;
            14'd10573: out = 12'hB47;
            14'd10574: out = 12'hB48;
            14'd10575: out = 12'hB48;
            14'd10576: out = 12'hB49;
            14'd10577: out = 12'hB49;
            14'd10578: out = 12'hB4A;
            14'd10579: out = 12'hB4A;
            14'd10580: out = 12'hB4B;
            14'd10581: out = 12'hB4B;
            14'd10582: out = 12'hB4C;
            14'd10583: out = 12'hB4C;
            14'd10584: out = 12'hB4D;
            14'd10585: out = 12'hB4D;
            14'd10586: out = 12'hB4E;
            14'd10587: out = 12'hB4E;
            14'd10588: out = 12'hB4F;
            14'd10589: out = 12'hB4F;
            14'd10590: out = 12'hB50;
            14'd10591: out = 12'hB50;
            14'd10592: out = 12'hB51;
            14'd10593: out = 12'hB51;
            14'd10594: out = 12'hB52;
            14'd10595: out = 12'hB52;
            14'd10596: out = 12'hB53;
            14'd10597: out = 12'hB53;
            14'd10598: out = 12'hB54;
            14'd10599: out = 12'hB54;
            14'd10600: out = 12'hB55;
            14'd10601: out = 12'hB55;
            14'd10602: out = 12'hB56;
            14'd10603: out = 12'hB56;
            14'd10604: out = 12'hB57;
            14'd10605: out = 12'hB57;
            14'd10606: out = 12'hB58;
            14'd10607: out = 12'hB58;
            14'd10608: out = 12'hB59;
            14'd10609: out = 12'hB59;
            14'd10610: out = 12'hB5A;
            14'd10611: out = 12'hB5A;
            14'd10612: out = 12'hB5B;
            14'd10613: out = 12'hB5B;
            14'd10614: out = 12'hB5C;
            14'd10615: out = 12'hB5C;
            14'd10616: out = 12'hB5D;
            14'd10617: out = 12'hB5D;
            14'd10618: out = 12'hB5E;
            14'd10619: out = 12'hB5E;
            14'd10620: out = 12'hB5F;
            14'd10621: out = 12'hB5F;
            14'd10622: out = 12'hB60;
            14'd10623: out = 12'hB60;
            14'd10624: out = 12'hB61;
            14'd10625: out = 12'hB61;
            14'd10626: out = 12'hB62;
            14'd10627: out = 12'hB62;
            14'd10628: out = 12'hB63;
            14'd10629: out = 12'hB63;
            14'd10630: out = 12'hB64;
            14'd10631: out = 12'hB64;
            14'd10632: out = 12'hB65;
            14'd10633: out = 12'hB65;
            14'd10634: out = 12'hB66;
            14'd10635: out = 12'hB66;
            14'd10636: out = 12'hB67;
            14'd10637: out = 12'hB67;
            14'd10638: out = 12'hB68;
            14'd10639: out = 12'hB68;
            14'd10640: out = 12'hB69;
            14'd10641: out = 12'hB69;
            14'd10642: out = 12'hB6A;
            14'd10643: out = 12'hB6A;
            14'd10644: out = 12'hB6B;
            14'd10645: out = 12'hB6B;
            14'd10646: out = 12'hB6C;
            14'd10647: out = 12'hB6C;
            14'd10648: out = 12'hB6D;
            14'd10649: out = 12'hB6D;
            14'd10650: out = 12'hB6E;
            default: out = 12'hB6F;
        endcase
    end
endmodule
