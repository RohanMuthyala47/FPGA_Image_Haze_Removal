module Transmission_Reciprocal_LUT (
    input      [9:0] in,  // Q0.10 input (unsigned, 0 to 0.65 range only)
    output reg [9:0] out  // Q2.8 reciprocal output (unsigned, 10-bit)
);

    always @(*) begin
        case(in)
            10'd  0: out = 10'h100;
            10'd  1: out = 10'h100;
            10'd  2: out = 10'h101;
            10'd  3: out = 10'h101;
            10'd  4: out = 10'h101;
            10'd  5: out = 10'h101;
            10'd  6: out = 10'h102;
            10'd  7: out = 10'h102;
            10'd  8: out = 10'h102;
            10'd  9: out = 10'h102;
            10'd 10: out = 10'h103;
            10'd 11: out = 10'h103;
            10'd 12: out = 10'h103;
            10'd 13: out = 10'h103;
            10'd 14: out = 10'h104;
            10'd 15: out = 10'h104;
            10'd 16: out = 10'h104;
            10'd 17: out = 10'h104;
            10'd 18: out = 10'h105;
            10'd 19: out = 10'h105;
            10'd 20: out = 10'h105;
            10'd 21: out = 10'h105;
            10'd 22: out = 10'h106;
            10'd 23: out = 10'h106;
            10'd 24: out = 10'h106;
            10'd 25: out = 10'h106;
            10'd 26: out = 10'h107;
            10'd 27: out = 10'h107;
            10'd 28: out = 10'h107;
            10'd 29: out = 10'h107;
            10'd 30: out = 10'h108;
            10'd 31: out = 10'h108;
            10'd 32: out = 10'h108;
            10'd 33: out = 10'h109;
            10'd 34: out = 10'h109;
            10'd 35: out = 10'h109;
            10'd 36: out = 10'h109;
            10'd 37: out = 10'h10A;
            10'd 38: out = 10'h10A;
            10'd 39: out = 10'h10A;
            10'd 40: out = 10'h10A;
            10'd 41: out = 10'h10B;
            10'd 42: out = 10'h10B;
            10'd 43: out = 10'h10B;
            10'd 44: out = 10'h10B;
            10'd 45: out = 10'h10C;
            10'd 46: out = 10'h10C;
            10'd 47: out = 10'h10C;
            10'd 48: out = 10'h10D;
            10'd 49: out = 10'h10D;
            10'd 50: out = 10'h10D;
            10'd 51: out = 10'h10D;
            10'd 52: out = 10'h10E;
            10'd 53: out = 10'h10E;
            10'd 54: out = 10'h10E;
            10'd 55: out = 10'h10F;
            10'd 56: out = 10'h10F;
            10'd 57: out = 10'h10F;
            10'd 58: out = 10'h10F;
            10'd 59: out = 10'h110;
            10'd 60: out = 10'h110;
            10'd 61: out = 10'h110;
            10'd 62: out = 10'h110;
            10'd 63: out = 10'h111;
            10'd 64: out = 10'h111;
            10'd 65: out = 10'h111;
            10'd 66: out = 10'h112;
            10'd 67: out = 10'h112;
            10'd 68: out = 10'h112;
            10'd 69: out = 10'h112;
            10'd 70: out = 10'h113;
            10'd 71: out = 10'h113;
            10'd 72: out = 10'h113;
            10'd 73: out = 10'h114;
            10'd 74: out = 10'h114;
            10'd 75: out = 10'h114;
            10'd 76: out = 10'h115;
            10'd 77: out = 10'h115;
            10'd 78: out = 10'h115;
            10'd 79: out = 10'h115;
            10'd 80: out = 10'h116;
            10'd 81: out = 10'h116;
            10'd 82: out = 10'h116;
            10'd 83: out = 10'h117;
            10'd 84: out = 10'h117;
            10'd 85: out = 10'h117;
            10'd 86: out = 10'h117;
            10'd 87: out = 10'h118;
            10'd 88: out = 10'h118;
            10'd 89: out = 10'h118;
            10'd 90: out = 10'h119;
            10'd 91: out = 10'h119;
            10'd 92: out = 10'h119;
            10'd 93: out = 10'h11A;
            10'd 94: out = 10'h11A;
            10'd 95: out = 10'h11A;
            10'd 96: out = 10'h11A;
            10'd 97: out = 10'h11B;
            10'd 98: out = 10'h11B;
            10'd 99: out = 10'h11B;
            10'd100: out = 10'h11C;
            10'd101: out = 10'h11C;
            10'd102: out = 10'h11C;
            10'd103: out = 10'h11D;
            10'd104: out = 10'h11D;
            10'd105: out = 10'h11D;
            10'd106: out = 10'h11E;
            10'd107: out = 10'h11E;
            10'd108: out = 10'h11E;
            10'd109: out = 10'h11E;
            10'd110: out = 10'h11F;
            10'd111: out = 10'h11F;
            10'd112: out = 10'h11F;
            10'd113: out = 10'h120;
            10'd114: out = 10'h120;
            10'd115: out = 10'h120;
            10'd116: out = 10'h121;
            10'd117: out = 10'h121;
            10'd118: out = 10'h121;
            10'd119: out = 10'h122;
            10'd120: out = 10'h122;
            10'd121: out = 10'h122;
            10'd122: out = 10'h123;
            10'd123: out = 10'h123;
            10'd124: out = 10'h123;
            10'd125: out = 10'h124;
            10'd126: out = 10'h124;
            10'd127: out = 10'h124;
            10'd128: out = 10'h125;
            10'd129: out = 10'h125;
            10'd130: out = 10'h125;
            10'd131: out = 10'h126;
            10'd132: out = 10'h126;
            10'd133: out = 10'h126;
            10'd134: out = 10'h127;
            10'd135: out = 10'h127;
            10'd136: out = 10'h127;
            10'd137: out = 10'h128;
            10'd138: out = 10'h128;
            10'd139: out = 10'h128;
            10'd140: out = 10'h129;
            10'd141: out = 10'h129;
            10'd142: out = 10'h129;
            10'd143: out = 10'h12A;
            10'd144: out = 10'h12A;
            10'd145: out = 10'h12A;
            10'd146: out = 10'h12B;
            10'd147: out = 10'h12B;
            10'd148: out = 10'h12B;
            10'd149: out = 10'h12C;
            10'd150: out = 10'h12C;
            10'd151: out = 10'h12C;
            10'd152: out = 10'h12D;
            10'd153: out = 10'h12D;
            10'd154: out = 10'h12D;
            10'd155: out = 10'h12E;
            10'd156: out = 10'h12E;
            10'd157: out = 10'h12E;
            10'd158: out = 10'h12F;
            10'd159: out = 10'h12F;
            10'd160: out = 10'h12F;
            10'd161: out = 10'h130;
            10'd162: out = 10'h130;
            10'd163: out = 10'h130;
            10'd164: out = 10'h131;
            10'd165: out = 10'h131;
            10'd166: out = 10'h132;
            10'd167: out = 10'h132;
            10'd168: out = 10'h132;
            10'd169: out = 10'h133;
            10'd170: out = 10'h133;
            10'd171: out = 10'h133;
            10'd172: out = 10'h134;
            10'd173: out = 10'h134;
            10'd174: out = 10'h134;
            10'd175: out = 10'h135;
            10'd176: out = 10'h135;
            10'd177: out = 10'h135;
            10'd178: out = 10'h136;
            10'd179: out = 10'h136;
            10'd180: out = 10'h137;
            10'd181: out = 10'h137;
            10'd182: out = 10'h137;
            10'd183: out = 10'h138;
            10'd184: out = 10'h138;
            10'd185: out = 10'h138;
            10'd186: out = 10'h139;
            10'd187: out = 10'h139;
            10'd188: out = 10'h13A;
            10'd189: out = 10'h13A;
            10'd190: out = 10'h13A;
            10'd191: out = 10'h13B;
            10'd192: out = 10'h13B;
            10'd193: out = 10'h13B;
            10'd194: out = 10'h13C;
            10'd195: out = 10'h13C;
            10'd196: out = 10'h13D;
            10'd197: out = 10'h13D;
            10'd198: out = 10'h13D;
            10'd199: out = 10'h13E;
            10'd200: out = 10'h13E;
            10'd201: out = 10'h13F;
            10'd202: out = 10'h13F;
            10'd203: out = 10'h13F;
            10'd204: out = 10'h140;
            10'd205: out = 10'h140;
            10'd206: out = 10'h140;
            10'd207: out = 10'h141;
            10'd208: out = 10'h141;
            10'd209: out = 10'h142;
            10'd210: out = 10'h142;
            10'd211: out = 10'h142;
            10'd212: out = 10'h143;
            10'd213: out = 10'h143;
            10'd214: out = 10'h144;
            10'd215: out = 10'h144;
            10'd216: out = 10'h144;
            10'd217: out = 10'h145;
            10'd218: out = 10'h145;
            10'd219: out = 10'h146;
            10'd220: out = 10'h146;
            10'd221: out = 10'h146;
            10'd222: out = 10'h147;
            10'd223: out = 10'h147;
            10'd224: out = 10'h148;
            10'd225: out = 10'h148;
            10'd226: out = 10'h149;
            10'd227: out = 10'h149;
            10'd228: out = 10'h149;
            10'd229: out = 10'h14A;
            10'd230: out = 10'h14A;
            10'd231: out = 10'h14B;
            10'd232: out = 10'h14B;
            10'd233: out = 10'h14B;
            10'd234: out = 10'h14C;
            10'd235: out = 10'h14C;
            10'd236: out = 10'h14D;
            10'd237: out = 10'h14D;
            10'd238: out = 10'h14E;
            10'd239: out = 10'h14E;
            10'd240: out = 10'h14E;
            10'd241: out = 10'h14F;
            10'd242: out = 10'h14F;
            10'd243: out = 10'h150;
            10'd244: out = 10'h150;
            10'd245: out = 10'h151;
            10'd246: out = 10'h151;
            10'd247: out = 10'h151;
            10'd248: out = 10'h152;
            10'd249: out = 10'h152;
            10'd250: out = 10'h153;
            10'd251: out = 10'h153;
            10'd252: out = 10'h154;
            10'd253: out = 10'h154;
            10'd254: out = 10'h154;
            10'd255: out = 10'h155;
            10'd256: out = 10'h155;
            10'd257: out = 10'h156;
            10'd258: out = 10'h156;
            10'd259: out = 10'h157;
            10'd260: out = 10'h157;
            10'd261: out = 10'h158;
            10'd262: out = 10'h158;
            10'd263: out = 10'h158;
            10'd264: out = 10'h159;
            10'd265: out = 10'h159;
            10'd266: out = 10'h15A;
            10'd267: out = 10'h15A;
            10'd268: out = 10'h15B;
            10'd269: out = 10'h15B;
            10'd270: out = 10'h15C;
            10'd271: out = 10'h15C;
            10'd272: out = 10'h15D;
            10'd273: out = 10'h15D;
            10'd274: out = 10'h15E;
            10'd275: out = 10'h15E;
            10'd276: out = 10'h15E;
            10'd277: out = 10'h15F;
            10'd278: out = 10'h15F;
            10'd279: out = 10'h160;
            10'd280: out = 10'h160;
            10'd281: out = 10'h161;
            10'd282: out = 10'h161;
            10'd283: out = 10'h162;
            10'd284: out = 10'h162;
            10'd285: out = 10'h163;
            10'd286: out = 10'h163;
            10'd287: out = 10'h164;
            10'd288: out = 10'h164;
            10'd289: out = 10'h165;
            10'd290: out = 10'h165;
            10'd291: out = 10'h166;
            10'd292: out = 10'h166;
            10'd293: out = 10'h167;
            10'd294: out = 10'h167;
            10'd295: out = 10'h168;
            10'd296: out = 10'h168;
            10'd297: out = 10'h169;
            10'd298: out = 10'h169;
            10'd299: out = 10'h16A;
            10'd300: out = 10'h16A;
            10'd301: out = 10'h16B;
            10'd302: out = 10'h16B;
            10'd303: out = 10'h16C;
            10'd304: out = 10'h16C;
            10'd305: out = 10'h16D;
            10'd306: out = 10'h16D;
            10'd307: out = 10'h16E;
            10'd308: out = 10'h16E;
            10'd309: out = 10'h16F;
            10'd310: out = 10'h16F;
            10'd311: out = 10'h170;
            10'd312: out = 10'h170;
            10'd313: out = 10'h171;
            10'd314: out = 10'h171;
            10'd315: out = 10'h172;
            10'd316: out = 10'h172;
            10'd317: out = 10'h173;
            10'd318: out = 10'h173;
            10'd319: out = 10'h174;
            10'd320: out = 10'h174;
            10'd321: out = 10'h175;
            10'd322: out = 10'h175;
            10'd323: out = 10'h176;
            10'd324: out = 10'h176;
            10'd325: out = 10'h177;
            10'd326: out = 10'h178;
            10'd327: out = 10'h178;
            10'd328: out = 10'h179;
            10'd329: out = 10'h179;
            10'd330: out = 10'h17A;
            10'd331: out = 10'h17A;
            10'd332: out = 10'h17B;
            10'd333: out = 10'h17B;
            10'd334: out = 10'h17C;
            10'd335: out = 10'h17C;
            10'd336: out = 10'h17D;
            10'd337: out = 10'h17E;
            10'd338: out = 10'h17E;
            10'd339: out = 10'h17F;
            10'd340: out = 10'h17F;
            10'd341: out = 10'h180;
            10'd342: out = 10'h180;
            10'd343: out = 10'h181;
            10'd344: out = 10'h182;
            10'd345: out = 10'h182;
            10'd346: out = 10'h183;
            10'd347: out = 10'h183;
            10'd348: out = 10'h184;
            10'd349: out = 10'h184;
            10'd350: out = 10'h185;
            10'd351: out = 10'h186;
            10'd352: out = 10'h186;
            10'd353: out = 10'h187;
            10'd354: out = 10'h187;
            10'd355: out = 10'h188;
            10'd356: out = 10'h188;
            10'd357: out = 10'h189;
            10'd358: out = 10'h18A;
            10'd359: out = 10'h18A;
            10'd360: out = 10'h18B;
            10'd361: out = 10'h18B;
            10'd362: out = 10'h18C;
            10'd363: out = 10'h18D;
            10'd364: out = 10'h18D;
            10'd365: out = 10'h18E;
            10'd366: out = 10'h18E;
            10'd367: out = 10'h18F;
            10'd368: out = 10'h190;
            10'd369: out = 10'h190;
            10'd370: out = 10'h191;
            10'd371: out = 10'h191;
            10'd372: out = 10'h192;
            10'd373: out = 10'h193;
            10'd374: out = 10'h193;
            10'd375: out = 10'h194;
            10'd376: out = 10'h195;
            10'd377: out = 10'h195;
            10'd378: out = 10'h196;
            10'd379: out = 10'h196;
            10'd380: out = 10'h197;
            10'd381: out = 10'h198;
            10'd382: out = 10'h198;
            10'd383: out = 10'h199;
            10'd384: out = 10'h19A;
            10'd385: out = 10'h19A;
            10'd386: out = 10'h19B;
            10'd387: out = 10'h19C;
            10'd388: out = 10'h19C;
            10'd389: out = 10'h19D;
            10'd390: out = 10'h19D;
            10'd391: out = 10'h19E;
            10'd392: out = 10'h19F;
            10'd393: out = 10'h19F;
            10'd394: out = 10'h1A0;
            10'd395: out = 10'h1A1;
            10'd396: out = 10'h1A1;
            10'd397: out = 10'h1A2;
            10'd398: out = 10'h1A3;
            10'd399: out = 10'h1A3;
            10'd400: out = 10'h1A4;
            10'd401: out = 10'h1A5;
            10'd402: out = 10'h1A5;
            10'd403: out = 10'h1A6;
            10'd404: out = 10'h1A7;
            10'd405: out = 10'h1A7;
            10'd406: out = 10'h1A8;
            10'd407: out = 10'h1A9;
            10'd408: out = 10'h1AA;
            10'd409: out = 10'h1AA;
            10'd410: out = 10'h1AB;
            10'd411: out = 10'h1AC;
            10'd412: out = 10'h1AC;
            10'd413: out = 10'h1AD;
            10'd414: out = 10'h1AE;
            10'd415: out = 10'h1AE;
            10'd416: out = 10'h1AF;
            10'd417: out = 10'h1B0;
            10'd418: out = 10'h1B1;
            10'd419: out = 10'h1B1;
            10'd420: out = 10'h1B2;
            10'd421: out = 10'h1B3;
            10'd422: out = 10'h1B3;
            10'd423: out = 10'h1B4;
            10'd424: out = 10'h1B5;
            10'd425: out = 10'h1B6;
            10'd426: out = 10'h1B6;
            10'd427: out = 10'h1B7;
            10'd428: out = 10'h1B8;
            10'd429: out = 10'h1B9;
            10'd430: out = 10'h1B9;
            10'd431: out = 10'h1BA;
            10'd432: out = 10'h1BB;
            10'd433: out = 10'h1BC;
            10'd434: out = 10'h1BC;
            10'd435: out = 10'h1BD;
            10'd436: out = 10'h1BE;
            10'd437: out = 10'h1BF;
            10'd438: out = 10'h1BF;
            10'd439: out = 10'h1C0;
            10'd440: out = 10'h1C1;
            10'd441: out = 10'h1C2;
            10'd442: out = 10'h1C2;
            10'd443: out = 10'h1C3;
            10'd444: out = 10'h1C4;
            10'd445: out = 10'h1C5;
            10'd446: out = 10'h1C6;
            10'd447: out = 10'h1C6;
            10'd448: out = 10'h1C7;
            10'd449: out = 10'h1C8;
            10'd450: out = 10'h1C9;
            10'd451: out = 10'h1C9;
            10'd452: out = 10'h1CA;
            10'd453: out = 10'h1CB;
            10'd454: out = 10'h1CC;
            10'd455: out = 10'h1CD;
            10'd456: out = 10'h1CE;
            10'd457: out = 10'h1CE;
            10'd458: out = 10'h1CF;
            10'd459: out = 10'h1D0;
            10'd460: out = 10'h1D1;
            10'd461: out = 10'h1D2;
            10'd462: out = 10'h1D2;
            10'd463: out = 10'h1D3;
            10'd464: out = 10'h1D4;
            10'd465: out = 10'h1D5;
            10'd466: out = 10'h1D6;
            10'd467: out = 10'h1D7;
            10'd468: out = 10'h1D7;
            10'd469: out = 10'h1D8;
            10'd470: out = 10'h1D9;
            10'd471: out = 10'h1DA;
            10'd472: out = 10'h1DB;
            10'd473: out = 10'h1DC;
            10'd474: out = 10'h1DD;
            10'd475: out = 10'h1DD;
            10'd476: out = 10'h1DE;
            10'd477: out = 10'h1DF;
            10'd478: out = 10'h1E0;
            10'd479: out = 10'h1E1;
            10'd480: out = 10'h1E2;
            10'd481: out = 10'h1E3;
            10'd482: out = 10'h1E4;
            10'd483: out = 10'h1E5;
            10'd484: out = 10'h1E5;
            10'd485: out = 10'h1E6;
            10'd486: out = 10'h1E7;
            10'd487: out = 10'h1E8;
            10'd488: out = 10'h1E9;
            10'd489: out = 10'h1EA;
            10'd490: out = 10'h1EB;
            10'd491: out = 10'h1EC;
            10'd492: out = 10'h1ED;
            10'd493: out = 10'h1EE;
            10'd494: out = 10'h1EF;
            10'd495: out = 10'h1F0;
            10'd496: out = 10'h1F0;
            10'd497: out = 10'h1F1;
            10'd498: out = 10'h1F2;
            10'd499: out = 10'h1F3;
            10'd500: out = 10'h1F4;
            10'd501: out = 10'h1F5;
            10'd502: out = 10'h1F6;
            10'd503: out = 10'h1F7;
            10'd504: out = 10'h1F8;
            10'd505: out = 10'h1F9;
            10'd506: out = 10'h1FA;
            10'd507: out = 10'h1FB;
            10'd508: out = 10'h1FC;
            10'd509: out = 10'h1FD;
            10'd510: out = 10'h1FE;
            10'd511: out = 10'h1FF;
            10'd512: out = 10'h200;
            10'd513: out = 10'h201;
            10'd514: out = 10'h202;
            10'd515: out = 10'h203;
            10'd516: out = 10'h204;
            10'd517: out = 10'h205;
            10'd518: out = 10'h206;
            10'd519: out = 10'h207;
            10'd520: out = 10'h208;
            10'd521: out = 10'h209;
            10'd522: out = 10'h20A;
            10'd523: out = 10'h20B;
            10'd524: out = 10'h20C;
            10'd525: out = 10'h20D;
            10'd526: out = 10'h20E;
            10'd527: out = 10'h20F;
            10'd528: out = 10'h211;
            10'd529: out = 10'h212;
            10'd530: out = 10'h213;
            10'd531: out = 10'h214;
            10'd532: out = 10'h215;
            10'd533: out = 10'h216;
            10'd534: out = 10'h217;
            10'd535: out = 10'h218;
            10'd536: out = 10'h219;
            10'd537: out = 10'h21A;
            10'd538: out = 10'h21B;
            10'd539: out = 10'h21D;
            10'd540: out = 10'h21E;
            10'd541: out = 10'h21F;
            10'd542: out = 10'h220;
            10'd543: out = 10'h221;
            10'd544: out = 10'h222;
            10'd545: out = 10'h223;
            10'd546: out = 10'h224;
            10'd547: out = 10'h226;
            10'd548: out = 10'h227;
            10'd549: out = 10'h228;
            10'd550: out = 10'h229;
            10'd551: out = 10'h22A;
            10'd552: out = 10'h22B;
            10'd553: out = 10'h22D;
            10'd554: out = 10'h22E;
            10'd555: out = 10'h22F;
            10'd556: out = 10'h230;
            10'd557: out = 10'h231;
            10'd558: out = 10'h233;
            10'd559: out = 10'h234;
            10'd560: out = 10'h235;
            10'd561: out = 10'h236;
            10'd562: out = 10'h237;
            10'd563: out = 10'h239;
            10'd564: out = 10'h23A;
            10'd565: out = 10'h23B;
            10'd566: out = 10'h23C;
            10'd567: out = 10'h23E;
            10'd568: out = 10'h23F;
            10'd569: out = 10'h240;
            10'd570: out = 10'h241;
            10'd571: out = 10'h243;
            10'd572: out = 10'h244;
            10'd573: out = 10'h245;
            10'd574: out = 10'h247;
            10'd575: out = 10'h248;
            10'd576: out = 10'h249;
            10'd577: out = 10'h24A;
            10'd578: out = 10'h24C;
            10'd579: out = 10'h24D;
            10'd580: out = 10'h24E;
            10'd581: out = 10'h250;
            10'd582: out = 10'h251;
            10'd583: out = 10'h252;
            10'd584: out = 10'h254;
            10'd585: out = 10'h255;
            10'd586: out = 10'h257;
            10'd587: out = 10'h258;
            10'd588: out = 10'h259;
            10'd589: out = 10'h25B;
            10'd590: out = 10'h25C;
            10'd591: out = 10'h25D;
            10'd592: out = 10'h25F;
            10'd593: out = 10'h260;
            10'd594: out = 10'h262;
            10'd595: out = 10'h263;
            10'd596: out = 10'h264;
            10'd597: out = 10'h266;
            10'd598: out = 10'h267;
            10'd599: out = 10'h269;
            10'd600: out = 10'h26A;
            10'd601: out = 10'h26C;
            10'd602: out = 10'h26D;
            10'd603: out = 10'h26F;
            10'd604: out = 10'h270;
            10'd605: out = 10'h272;
            10'd606: out = 10'h273;
            10'd607: out = 10'h275;
            10'd608: out = 10'h276;
            10'd609: out = 10'h278;
            10'd610: out = 10'h279;
            10'd611: out = 10'h27B;
            10'd612: out = 10'h27C;
            10'd613: out = 10'h27E;
            10'd614: out = 10'h27F;
            10'd615: out = 10'h281;
            10'd616: out = 10'h283;
            10'd617: out = 10'h284;
            10'd618: out = 10'h286;
            10'd619: out = 10'h287;
            10'd620: out = 10'h289;
            10'd621: out = 10'h28A;
            10'd622: out = 10'h28C;
            10'd623: out = 10'h28E;
            10'd624: out = 10'h28F;
            10'd625: out = 10'h291;
            10'd626: out = 10'h293;
            10'd627: out = 10'h294;
            10'd628: out = 10'h296;
            10'd629: out = 10'h298;
            10'd630: out = 10'h299;
            10'd631: out = 10'h29B;
            10'd632: out = 10'h29D;
            10'd633: out = 10'h29E;
            10'd634: out = 10'h2A0;
            10'd635: out = 10'h2A2;
            10'd636: out = 10'h2A4;
            10'd637: out = 10'h2A5;
            10'd638: out = 10'h2A7;
            10'd639: out = 10'h2A9;
            10'd640: out = 10'h2AB;
            10'd641: out = 10'h2AC;
            10'd642: out = 10'h2AE;
            10'd643: out = 10'h2B0;
            10'd644: out = 10'h2B2;
            10'd645: out = 10'h2B4;
            10'd646: out = 10'h2B6;
            10'd647: out = 10'h2B7;
            10'd648: out = 10'h2B9;
            10'd649: out = 10'h2BB;
            10'd650: out = 10'h2BD;
            10'd651: out = 10'h2BF;
            10'd652: out = 10'h2C1;
            10'd653: out = 10'h2C3;
            10'd654: out = 10'h2C4;
            10'd655: out = 10'h2C6;
            10'd656: out = 10'h2C8;
            10'd657: out = 10'h2CA;
            10'd658: out = 10'h2CC;
            10'd659: out = 10'h2CE;
            10'd660: out = 10'h2D0;
            10'd661: out = 10'h2D2;
            10'd662: out = 10'h2D4;
            10'd663: out = 10'h2D6;
            10'd664: out = 10'h2D8;
            10'd665: out = 10'h2DA;
            10'd666: out = 10'h2DC;
            default: out = 10'h2DE;
        endcase
    end
    
endmodule
