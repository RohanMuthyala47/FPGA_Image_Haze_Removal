module Atmospheric_Light_Reciprocal_LUT (
    input  [7:0] in,
    output reg [9:0] out
);

    always @(*) begin
        casez (in)
            8'd  1: out = 10'd 960;  // 0.9375/1 ≈ 0.93750000
            8'd  2: out = 10'd 480;  // 0.9375/2 ≈ 0.46875000
            8'd  3: out = 10'd 320;  // 0.9375/3 ≈ 0.31250000
            8'd  4: out = 10'd 240;  // 0.9375/4 ≈ 0.23437500
            8'd  5: out = 10'd 192;  // 0.9375/5 ≈ 0.18750000
            8'd  6: out = 10'd 160;  // 0.9375/6 ≈ 0.15625000
            8'd  7: out = 10'd 137;  // 0.9375/7 ≈ 0.13392857
            8'd  8: out = 10'd 120;  // 0.9375/8 ≈ 0.11718750
            8'd  9: out = 10'd 107;  // 0.9375/9 ≈ 0.10416667
            8'd 10: out = 10'd  96;  // 0.9375/10 ≈ 0.09375000
            8'd 11: out = 10'd  87;  // 0.9375/11 ≈ 0.08522727
            8'd 12: out = 10'd  80;  // 0.9375/12 ≈ 0.07812500
            8'd 13: out = 10'd  74;  // 0.9375/13 ≈ 0.07211538
            8'd 14: out = 10'd  69;  // 0.9375/14 ≈ 0.06696429
            8'd 15: out = 10'd  64;  // 0.9375/15 ≈ 0.06250000
            8'd 16: out = 10'd  60;  // 0.9375/16 ≈ 0.05859375
            8'd 17: out = 10'd  56;  // 0.9375/17 ≈ 0.05514706
            8'd 18: out = 10'd  53;  // 0.9375/18 ≈ 0.05208333
            8'd 19: out = 10'd  51;  // 0.9375/19 ≈ 0.04934211
            8'd 20: out = 10'd  48;  // 0.9375/20 ≈ 0.04687500
            8'd 21: out = 10'd  46;  // 0.9375/21 ≈ 0.04464286
            8'd 22: out = 10'd  44;  // 0.9375/22 ≈ 0.04261364
            8'd 23: out = 10'd  42;  // 0.9375/23 ≈ 0.04076087
            8'd 24: out = 10'd  40;  // 0.9375/24 ≈ 0.03906250
            8'd 25: out = 10'd  38;  // 0.9375/25 ≈ 0.03750000
            8'd 26: out = 10'd  37;  // 0.9375/26 ≈ 0.03605769
            8'd 27: out = 10'd  36;  // 0.9375/27 ≈ 0.03472222
            8'd 28: out = 10'd  34;  // 0.9375/28 ≈ 0.03348214
            8'd 29: out = 10'd  33;  // 0.9375/29 ≈ 0.03232759
            8'd 30: out = 10'd  32;  // 0.9375/30 ≈ 0.03125000
            8'd 31: out = 10'd  31;  // 0.9375/31 ≈ 0.03024194
            8'd 32: out = 10'd  30;  // 0.9375/32 ≈ 0.02929688
            8'd 33: out = 10'd  29;  // 0.9375/33 ≈ 0.02840909
            8'd 34: out = 10'd  28;  // 0.9375/34 ≈ 0.02757353
            8'd 35: out = 10'd  27;  // 0.9375/35 ≈ 0.02678571
            8'd 36: out = 10'd  27;  // 0.9375/36 ≈ 0.02604167
            8'd 37: out = 10'd  26;  // 0.9375/37 ≈ 0.02533784
            8'd 38: out = 10'd  25;  // 0.9375/38 ≈ 0.02467105
            8'd 39: out = 10'd  25;  // 0.9375/39 ≈ 0.02403846
            8'd 40: out = 10'd  24;  // 0.9375/40 ≈ 0.02343750
            8'd 41: out = 10'd  23;  // 0.9375/41 ≈ 0.02286585
            8'd 42: out = 10'd  23;  // 0.9375/42 ≈ 0.02232143
            8'd 43: out = 10'd  22;  // 0.9375/43 ≈ 0.02180233
            8'd 44: out = 10'd  22;  // 0.9375/44 ≈ 0.02130682
            8'd 45: out = 10'd  21;  // 0.9375/45 ≈ 0.02083333
            8'd 46: out = 10'd  21;  // 0.9375/46 ≈ 0.02038043
            8'd 47: out = 10'd  20;  // 0.9375/47 ≈ 0.01994681
            8'd 48: out = 10'd  20;  // 0.9375/48 ≈ 0.01953125
            8'd 49: out = 10'd  20;  // 0.9375/49 ≈ 0.01913265
            8'd 50: out = 10'd  19;  // 0.9375/50 ≈ 0.01875000
            8'd 51: out = 10'd  19;  // 0.9375/51 ≈ 0.01838235
            8'd 52: out = 10'd  18;  // 0.9375/52 ≈ 0.01802885
            8'd 53: out = 10'd  18;  // 0.9375/53 ≈ 0.01768868
            8'd 54: out = 10'd  18;  // 0.9375/54 ≈ 0.01736111
            8'd 55: out = 10'd  17;  // 0.9375/55 ≈ 0.01704545
            8'd 56: out = 10'd  17;  // 0.9375/56 ≈ 0.01674107
            8'd 57: out = 10'd  17;  // 0.9375/57 ≈ 0.01644737
            8'd 58: out = 10'd  17;  // 0.9375/58 ≈ 0.01616379
            8'd 59: out = 10'd  16;  // 0.9375/59 ≈ 0.01588983
            8'd 60: out = 10'd  16;  // 0.9375/60 ≈ 0.01562500
            8'd 61: out = 10'd  16;  // 0.9375/61 ≈ 0.01536885
            8'd 62: out = 10'd  15;  // 0.9375/62 ≈ 0.01512097
            8'd 63: out = 10'd  15;  // 0.9375/63 ≈ 0.01488095
            8'd 64: out = 10'd  15;  // 0.9375/64 ≈ 0.01464844
            8'd 65: out = 10'd  15;  // 0.9375/65 ≈ 0.01442308
            8'd 66: out = 10'd  15;  // 0.9375/66 ≈ 0.01420455
            8'd 67: out = 10'd  14;  // 0.9375/67 ≈ 0.01399254
            8'd 68: out = 10'd  14;  // 0.9375/68 ≈ 0.01378676
            8'd 69: out = 10'd  14;  // 0.9375/69 ≈ 0.01358696
            8'd 70: out = 10'd  14;  // 0.9375/70 ≈ 0.01339286
            8'd 71: out = 10'd  14;  // 0.9375/71 ≈ 0.01320423
            8'd 72: out = 10'd  13;  // 0.9375/72 ≈ 0.01302083
            8'd 73: out = 10'd  13;  // 0.9375/73 ≈ 0.01284247
            8'd 74: out = 10'd  13;  // 0.9375/74 ≈ 0.01266892
            8'd 75: out = 10'd  13;  // 0.9375/75 ≈ 0.01250000
            8'd 76: out = 10'd  13;  // 0.9375/76 ≈ 0.01233553
            8'd 77: out = 10'd  12;  // 0.9375/77 ≈ 0.01217532
            8'd 78: out = 10'd  12;  // 0.9375/78 ≈ 0.01201923
            8'd 79: out = 10'd  12;  // 0.9375/79 ≈ 0.01186709
            8'd 80: out = 10'd  12;  // 0.9375/80 ≈ 0.01171875
            8'd 81: out = 10'd  12;  // 0.9375/81 ≈ 0.01157407
            8'd 82: out = 10'd  12;  // 0.9375/82 ≈ 0.01143293
            8'd 83: out = 10'd  12;  // 0.9375/83 ≈ 0.01129518
            8'd 84: out = 10'd  11;  // 0.9375/84 ≈ 0.01116071
            8'd 85: out = 10'd  11;  // 0.9375/85 ≈ 0.01102941
            8'd 86: out = 10'd  11;  // 0.9375/86 ≈ 0.01090116
            8'd 87: out = 10'd  11;  // 0.9375/87 ≈ 0.01077586
            8'd 88: out = 10'd  11;  // 0.9375/88 ≈ 0.01065341
            8'd 89: out = 10'd  11;  // 0.9375/89 ≈ 0.01053371
            8'd 90: out = 10'd  11;  // 0.9375/90 ≈ 0.01041667
            8'd 91: out = 10'd  11;  // 0.9375/91 ≈ 0.01030220
            8'd 92: out = 10'd  10;  // 0.9375/92 ≈ 0.01019022
            8'd 93: out = 10'd  10;  // 0.9375/93 ≈ 0.01008065
            8'd 94: out = 10'd  10;  // 0.9375/94 ≈ 0.00997340
            8'd 95: out = 10'd  10;  // 0.9375/95 ≈ 0.00986842
            8'd 96: out = 10'd  10;  // 0.9375/96 ≈ 0.00976562
            8'd 97: out = 10'd  10;  // 0.9375/97 ≈ 0.00966495
            8'd 98: out = 10'd  10;  // 0.9375/98 ≈ 0.00956633
            8'd 99: out = 10'd  10;  // 0.9375/99 ≈ 0.00946970
            8'd100: out = 10'd  10;  // 0.9375/100 ≈ 0.00937500
            8'd101: out = 10'd  10;  // 0.9375/101 ≈ 0.00928218
            8'd102: out = 10'd   9;  // 0.9375/102 ≈ 0.00919118
            8'd103: out = 10'd   9;  // 0.9375/103 ≈ 0.00910194
            8'd104: out = 10'd   9;  // 0.9375/104 ≈ 0.00901442
            8'd105: out = 10'd   9;  // 0.9375/105 ≈ 0.00892857
            8'd106: out = 10'd   9;  // 0.9375/106 ≈ 0.00884434
            8'd107: out = 10'd   9;  // 0.9375/107 ≈ 0.00876168
            8'd108: out = 10'd   9;  // 0.9375/108 ≈ 0.00868056
            8'd109: out = 10'd   9;  // 0.9375/109 ≈ 0.00860092
            8'd110: out = 10'd   9;  // 0.9375/110 ≈ 0.00852273
            8'd111: out = 10'd   9;  // 0.9375/111 ≈ 0.00844595
            8'd112: out = 10'd   9;  // 0.9375/112 ≈ 0.00837054
            8'd113: out = 10'd   8;  // 0.9375/113 ≈ 0.00829646
            8'd114: out = 10'd   8;  // 0.9375/114 ≈ 0.00822368
            8'd115: out = 10'd   8;  // 0.9375/115 ≈ 0.00815217
            8'd116: out = 10'd   8;  // 0.9375/116 ≈ 0.00808190
            8'd117: out = 10'd   8;  // 0.9375/117 ≈ 0.00801282
            8'd118: out = 10'd   8;  // 0.9375/118 ≈ 0.00794492
            8'd119: out = 10'd   8;  // 0.9375/119 ≈ 0.00787815
            8'd120: out = 10'd   8;  // 0.9375/120 ≈ 0.00781250
            8'd121: out = 10'd   8;  // 0.9375/121 ≈ 0.00774793
            8'd122: out = 10'd   8;  // 0.9375/122 ≈ 0.00768443
            8'd123: out = 10'd   8;  // 0.9375/123 ≈ 0.00762195
            8'd124: out = 10'd   8;  // 0.9375/124 ≈ 0.00756048
            8'd125: out = 10'd   8;  // 0.9375/125 ≈ 0.00750000
            8'd126: out = 10'd   8;  // 0.9375/126 ≈ 0.00744048
            8'd127: out = 10'd   8;  // 0.9375/127 ≈ 0.00738189
            8'd128: out = 10'd   8;  // 0.9375/128 ≈ 0.00732422
            8'd129: out = 10'd   7;  // 0.9375/129 ≈ 0.00726744
            8'd130: out = 10'd   7;  // 0.9375/130 ≈ 0.00721154
            8'd131: out = 10'd   7;  // 0.9375/131 ≈ 0.00715649
            8'd132: out = 10'd   7;  // 0.9375/132 ≈ 0.00710227
            8'd133: out = 10'd   7;  // 0.9375/133 ≈ 0.00704887
            8'd134: out = 10'd   7;  // 0.9375/134 ≈ 0.00699627
            8'd135: out = 10'd   7;  // 0.9375/135 ≈ 0.00694444
            8'd136: out = 10'd   7;  // 0.9375/136 ≈ 0.00689338
            8'd137: out = 10'd   7;  // 0.9375/137 ≈ 0.00684307
            8'd138: out = 10'd   7;  // 0.9375/138 ≈ 0.00679348
            8'd139: out = 10'd   7;  // 0.9375/139 ≈ 0.00674460
            8'd140: out = 10'd   7;  // 0.9375/140 ≈ 0.00669643
            8'd141: out = 10'd   7;  // 0.9375/141 ≈ 0.00664894
            8'd142: out = 10'd   7;  // 0.9375/142 ≈ 0.00660211
            8'd143: out = 10'd   7;  // 0.9375/143 ≈ 0.00655594
            8'd144: out = 10'd   7;  // 0.9375/144 ≈ 0.00651042
            8'd145: out = 10'd   7;  // 0.9375/145 ≈ 0.00646552
            8'd146: out = 10'd   7;  // 0.9375/146 ≈ 0.00642123
            8'd147: out = 10'd   7;  // 0.9375/147 ≈ 0.00637755
            8'd148: out = 10'd   6;  // 0.9375/148 ≈ 0.00633446
            8'd149: out = 10'd   6;  // 0.9375/149 ≈ 0.00629195
            8'd150: out = 10'd   6;  // 0.9375/150 ≈ 0.00625000
            8'd151: out = 10'd   6;  // 0.9375/151 ≈ 0.00620861
            8'd152: out = 10'd   6;  // 0.9375/152 ≈ 0.00616776
            8'd153: out = 10'd   6;  // 0.9375/153 ≈ 0.00612745
            8'd154: out = 10'd   6;  // 0.9375/154 ≈ 0.00608766
            8'd155: out = 10'd   6;  // 0.9375/155 ≈ 0.00604839
            8'd156: out = 10'd   6;  // 0.9375/156 ≈ 0.00600962
            8'd157: out = 10'd   6;  // 0.9375/157 ≈ 0.00597134
            8'd158: out = 10'd   6;  // 0.9375/158 ≈ 0.00593354
            8'd159: out = 10'd   6;  // 0.9375/159 ≈ 0.00589623
            8'd160: out = 10'd   6;  // 0.9375/160 ≈ 0.00585938
            8'd161: out = 10'd   6;  // 0.9375/161 ≈ 0.00582298
            8'd162: out = 10'd   6;  // 0.9375/162 ≈ 0.00578704
            8'd163: out = 10'd   6;  // 0.9375/163 ≈ 0.00575153
            8'd164: out = 10'd   6;  // 0.9375/164 ≈ 0.00571646
            8'd165: out = 10'd   6;  // 0.9375/165 ≈ 0.00568182
            8'd166: out = 10'd   6;  // 0.9375/166 ≈ 0.00564759
            8'd167: out = 10'd   6;  // 0.9375/167 ≈ 0.00561377
            8'd168: out = 10'd   6;  // 0.9375/168 ≈ 0.00558036
            8'd169: out = 10'd   6;  // 0.9375/169 ≈ 0.00554734
            8'd170: out = 10'd   6;  // 0.9375/170 ≈ 0.00551471
            8'd171: out = 10'd   6;  // 0.9375/171 ≈ 0.00548246
            8'd172: out = 10'd   6;  // 0.9375/172 ≈ 0.00545058
            8'd173: out = 10'd   6;  // 0.9375/173 ≈ 0.00541908
            8'd174: out = 10'd   6;  // 0.9375/174 ≈ 0.00538793
            8'd175: out = 10'd   5;  // 0.9375/175 ≈ 0.00535714
            8'd176: out = 10'd   5;  // 0.9375/176 ≈ 0.00532670
            8'd177: out = 10'd   5;  // 0.9375/177 ≈ 0.00529661
            8'd178: out = 10'd   5;  // 0.9375/178 ≈ 0.00526685
            8'd179: out = 10'd   5;  // 0.9375/179 ≈ 0.00523743
            8'd180: out = 10'd   5;  // 0.9375/180 ≈ 0.00520833
            8'd181: out = 10'd   5;  // 0.9375/181 ≈ 0.00517956
            8'd182: out = 10'd   5;  // 0.9375/182 ≈ 0.00515110
            8'd183: out = 10'd   5;  // 0.9375/183 ≈ 0.00512295
            8'd184: out = 10'd   5;  // 0.9375/184 ≈ 0.00509511
            8'd185: out = 10'd   5;  // 0.9375/185 ≈ 0.00506757
            8'd186: out = 10'd   5;  // 0.9375/186 ≈ 0.00504032
            8'd187: out = 10'd   5;  // 0.9375/187 ≈ 0.00501337
            8'd188: out = 10'd   5;  // 0.9375/188 ≈ 0.00498670
            8'd189: out = 10'd   5;  // 0.9375/189 ≈ 0.00496032
            8'd190: out = 10'd   5;  // 0.9375/190 ≈ 0.00493421
            8'd191: out = 10'd   5;  // 0.9375/191 ≈ 0.00490838
            8'd192: out = 10'd   5;  // 0.9375/192 ≈ 0.00488281
            8'd193: out = 10'd   5;  // 0.9375/193 ≈ 0.00485751
            8'd194: out = 10'd   5;  // 0.9375/194 ≈ 0.00483247
            8'd195: out = 10'd   5;  // 0.9375/195 ≈ 0.00480769
            8'd196: out = 10'd   5;  // 0.9375/196 ≈ 0.00478316
            8'd197: out = 10'd   5;  // 0.9375/197 ≈ 0.00475888
            8'd198: out = 10'd   5;  // 0.9375/198 ≈ 0.00473485
            8'd199: out = 10'd   5;  // 0.9375/199 ≈ 0.00471106
            8'd200: out = 10'd   5;  // 0.9375/200 ≈ 0.00468750
            8'd201: out = 10'd   5;  // 0.9375/201 ≈ 0.00466418
            8'd202: out = 10'd   5;  // 0.9375/202 ≈ 0.00464109
            8'd203: out = 10'd   5;  // 0.9375/203 ≈ 0.00461823
            8'd204: out = 10'd   5;  // 0.9375/204 ≈ 0.00459559
            8'd205: out = 10'd   5;  // 0.9375/205 ≈ 0.00457317
            8'd206: out = 10'd   5;  // 0.9375/206 ≈ 0.00455097
            8'd207: out = 10'd   5;  // 0.9375/207 ≈ 0.00452899
            8'd208: out = 10'd   5;  // 0.9375/208 ≈ 0.00450721
            8'd209: out = 10'd   5;  // 0.9375/209 ≈ 0.00448565
            8'd210: out = 10'd   5;  // 0.9375/210 ≈ 0.00446429
            8'd211: out = 10'd   5;  // 0.9375/211 ≈ 0.00444313
            8'd212: out = 10'd   5;  // 0.9375/212 ≈ 0.00442217
            8'd213: out = 10'd   5;  // 0.9375/213 ≈ 0.00440141
            8'd214: out = 10'd   4;  // 0.9375/214 ≈ 0.00438084
            8'd215: out = 10'd   4;  // 0.9375/215 ≈ 0.00436047
            8'd216: out = 10'd   4;  // 0.9375/216 ≈ 0.00434028
            8'd217: out = 10'd   4;  // 0.9375/217 ≈ 0.00432028
            8'd218: out = 10'd   4;  // 0.9375/218 ≈ 0.00430046
            8'd219: out = 10'd   4;  // 0.9375/219 ≈ 0.00428082
            8'd220: out = 10'd   4;  // 0.9375/220 ≈ 0.00426136
            8'd221: out = 10'd   4;  // 0.9375/221 ≈ 0.00424208
            8'd222: out = 10'd   4;  // 0.9375/222 ≈ 0.00422297
            8'd223: out = 10'd   4;  // 0.9375/223 ≈ 0.00420404
            8'd224: out = 10'd   4;  // 0.9375/224 ≈ 0.00418527
            8'd225: out = 10'd   4;  // 0.9375/225 ≈ 0.00416667
            8'd226: out = 10'd   4;  // 0.9375/226 ≈ 0.00414823
            8'd227: out = 10'd   4;  // 0.9375/227 ≈ 0.00412996
            8'd228: out = 10'd   4;  // 0.9375/228 ≈ 0.00411184
            8'd229: out = 10'd   4;  // 0.9375/229 ≈ 0.00409389
            8'd230: out = 10'd   4;  // 0.9375/230 ≈ 0.00407609
            8'd231: out = 10'd   4;  // 0.9375/231 ≈ 0.00405844
            8'd232: out = 10'd   4;  // 0.9375/232 ≈ 0.00404095
            8'd233: out = 10'd   4;  // 0.9375/233 ≈ 0.00402361
            8'd234: out = 10'd   4;  // 0.9375/234 ≈ 0.00400641
            8'd235: out = 10'd   4;  // 0.9375/235 ≈ 0.00398936
            8'd236: out = 10'd   4;  // 0.9375/236 ≈ 0.00397246
            8'd237: out = 10'd   4;  // 0.9375/237 ≈ 0.00395570
            8'd238: out = 10'd   4;  // 0.9375/238 ≈ 0.00393908
            8'd239: out = 10'd   4;  // 0.9375/239 ≈ 0.00392259
            8'd240: out = 10'd   4;  // 0.9375/240 ≈ 0.00390625
            8'd241: out = 10'd   4;  // 0.9375/241 ≈ 0.00389004
            8'd242: out = 10'd   4;  // 0.9375/242 ≈ 0.00387397
            8'd243: out = 10'd   4;  // 0.9375/243 ≈ 0.00385802
            8'd244: out = 10'd   4;  // 0.9375/244 ≈ 0.00384221
            8'd245: out = 10'd   4;  // 0.9375/245 ≈ 0.00382653
            8'd246: out = 10'd   4;  // 0.9375/246 ≈ 0.00381098
            8'd247: out = 10'd   4;  // 0.9375/247 ≈ 0.00379555
            8'd248: out = 10'd   4;  // 0.9375/248 ≈ 0.00378024
            8'd249: out = 10'd   4;  // 0.9375/249 ≈ 0.00376506
            8'd250: out = 10'd   4;  // 0.9375/250 ≈ 0.00375000
            8'd251: out = 10'd   4;  // 0.9375/251 ≈ 0.00373506
            8'd252: out = 10'd   4;  // 0.9375/252 ≈ 0.00372024
            8'd253: out = 10'd   4;  // 0.9375/253 ≈ 0.00370553
            8'd254: out = 10'd   4;  // 0.9375/254 ≈ 0.00369094
            8'd255: out = 10'd   4;  // 0.9375/255 ≈ 0.00367647
            default: out = 10'd1023; // default case
        endcase
    end

endmodule
