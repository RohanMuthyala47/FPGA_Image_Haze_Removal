module Atmospheric_Light_Reciprocal_LUT (
    input      [7:0] in,
    output reg [13:0] out
);

    always @(*) begin
        case (in)
            8'd  1: out = 14'd16383;  // 1/1 ? 1.00000000
            8'd  2: out = 14'd 8192;  // 1/2 ? 0.50000000
            8'd  3: out = 14'd 5461;  // 1/3 ? 0.33333333
            8'd  4: out = 14'd 4096;  // 1/4 ? 0.25000000
            8'd  5: out = 14'd 3277;  // 1/5 ? 0.20000000
            8'd  6: out = 14'd 2731;  // 1/6 ? 0.16666667
            8'd  7: out = 14'd 2341;  // 1/7 ? 0.14285714
            8'd  8: out = 14'd 2048;  // 1/8 ? 0.12500000
            8'd  9: out = 14'd 1820;  // 1/9 ? 0.11111111
            8'd 10: out = 14'd 1638;  // 1/10 ? 0.10000000
            8'd 11: out = 14'd 1489;  // 1/11 ? 0.09090909
            8'd 12: out = 14'd 1365;  // 1/12 ? 0.08333333
            8'd 13: out = 14'd 1260;  // 1/13 ? 0.07692308
            8'd 14: out = 14'd 1170;  // 1/14 ? 0.07142857
            8'd 15: out = 14'd 1092;  // 1/15 ? 0.06666667
            8'd 16: out = 14'd 1024;  // 1/16 ? 0.06250000
            8'd 17: out = 14'd  964;  // 1/17 ? 0.05882353
            8'd 18: out = 14'd  910;  // 1/18 ? 0.05555556
            8'd 19: out = 14'd  862;  // 1/19 ? 0.05263158
            8'd 20: out = 14'd  819;  // 1/20 ? 0.05000000
            8'd 21: out = 14'd  780;  // 1/21 ? 0.04761905
            8'd 22: out = 14'd  745;  // 1/22 ? 0.04545455
            8'd 23: out = 14'd  712;  // 1/23 ? 0.04347826
            8'd 24: out = 14'd  683;  // 1/24 ? 0.04166667
            8'd 25: out = 14'd  655;  // 1/25 ? 0.04000000
            8'd 26: out = 14'd  630;  // 1/26 ? 0.03846154
            8'd 27: out = 14'd  607;  // 1/27 ? 0.03703704
            8'd 28: out = 14'd  585;  // 1/28 ? 0.03571429
            8'd 29: out = 14'd  565;  // 1/29 ? 0.03448276
            8'd 30: out = 14'd  546;  // 1/30 ? 0.03333333
            8'd 31: out = 14'd  529;  // 1/31 ? 0.03225806
            8'd 32: out = 14'd  512;  // 1/32 ? 0.03125000
            8'd 33: out = 14'd  496;  // 1/33 ? 0.03030303
            8'd 34: out = 14'd  482;  // 1/34 ? 0.02941176
            8'd 35: out = 14'd  468;  // 1/35 ? 0.02857143
            8'd 36: out = 14'd  455;  // 1/36 ? 0.02777778
            8'd 37: out = 14'd  443;  // 1/37 ? 0.02702703
            8'd 38: out = 14'd  431;  // 1/38 ? 0.02631579
            8'd 39: out = 14'd  420;  // 1/39 ? 0.02564103
            8'd 40: out = 14'd  410;  // 1/40 ? 0.02500000
            8'd 41: out = 14'd  400;  // 1/41 ? 0.02439024
            8'd 42: out = 14'd  390;  // 1/42 ? 0.02380952
            8'd 43: out = 14'd  381;  // 1/43 ? 0.02325581
            8'd 44: out = 14'd  372;  // 1/44 ? 0.02272727
            8'd 45: out = 14'd  364;  // 1/45 ? 0.02222222
            8'd 46: out = 14'd  356;  // 1/46 ? 0.02173913
            8'd 47: out = 14'd  349;  // 1/47 ? 0.02127660
            8'd 48: out = 14'd  341;  // 1/48 ? 0.02083333
            8'd 49: out = 14'd  334;  // 1/49 ? 0.02040816
            8'd 50: out = 14'd  328;  // 1/50 ? 0.02000000
            8'd 51: out = 14'd  321;  // 1/51 ? 0.01960784
            8'd 52: out = 14'd  315;  // 1/52 ? 0.01923077
            8'd 53: out = 14'd  309;  // 1/53 ? 0.01886792
            8'd 54: out = 14'd  303;  // 1/54 ? 0.01851852
            8'd 55: out = 14'd  298;  // 1/55 ? 0.01818182
            8'd 56: out = 14'd  293;  // 1/56 ? 0.01785714
            8'd 57: out = 14'd  287;  // 1/57 ? 0.01754386
            8'd 58: out = 14'd  282;  // 1/58 ? 0.01724138
            8'd 59: out = 14'd  278;  // 1/59 ? 0.01694915
            8'd 60: out = 14'd  273;  // 1/60 ? 0.01666667
            8'd 61: out = 14'd  269;  // 1/61 ? 0.01639344
            8'd 62: out = 14'd  264;  // 1/62 ? 0.01612903
            8'd 63: out = 14'd  260;  // 1/63 ? 0.01587302
            8'd 64: out = 14'd  256;  // 1/64 ? 0.01562500
            8'd 65: out = 14'd  252;  // 1/65 ? 0.01538462
            8'd 66: out = 14'd  248;  // 1/66 ? 0.01515152
            8'd 67: out = 14'd  245;  // 1/67 ? 0.01492537
            8'd 68: out = 14'd  241;  // 1/68 ? 0.01470588
            8'd 69: out = 14'd  237;  // 1/69 ? 0.01449275
            8'd 70: out = 14'd  234;  // 1/70 ? 0.01428571
            8'd 71: out = 14'd  231;  // 1/71 ? 0.01408451
            8'd 72: out = 14'd  228;  // 1/72 ? 0.01388889
            8'd 73: out = 14'd  224;  // 1/73 ? 0.01369863
            8'd 74: out = 14'd  221;  // 1/74 ? 0.01351351
            8'd 75: out = 14'd  218;  // 1/75 ? 0.01333333
            8'd 76: out = 14'd  216;  // 1/76 ? 0.01315789
            8'd 77: out = 14'd  213;  // 1/77 ? 0.01298701
            8'd 78: out = 14'd  210;  // 1/78 ? 0.01282051
            8'd 79: out = 14'd  207;  // 1/79 ? 0.01265823
            8'd 80: out = 14'd  205;  // 1/80 ? 0.01250000
            8'd 81: out = 14'd  202;  // 1/81 ? 0.01234568
            8'd 82: out = 14'd  200;  // 1/82 ? 0.01219512
            8'd 83: out = 14'd  197;  // 1/83 ? 0.01204819
            8'd 84: out = 14'd  195;  // 1/84 ? 0.01190476
            8'd 85: out = 14'd  193;  // 1/85 ? 0.01176471
            8'd 86: out = 14'd  191;  // 1/86 ? 0.01162791
            8'd 87: out = 14'd  188;  // 1/87 ? 0.01149425
            8'd 88: out = 14'd  186;  // 1/88 ? 0.01136364
            8'd 89: out = 14'd  184;  // 1/89 ? 0.01123596
            8'd 90: out = 14'd  182;  // 1/90 ? 0.01111111
            8'd 91: out = 14'd  180;  // 1/91 ? 0.01098901
            8'd 92: out = 14'd  178;  // 1/92 ? 0.01086957
            8'd 93: out = 14'd  176;  // 1/93 ? 0.01075269
            8'd 94: out = 14'd  174;  // 1/94 ? 0.01063830
            8'd 95: out = 14'd  172;  // 1/95 ? 0.01052632
            8'd 96: out = 14'd  171;  // 1/96 ? 0.01041667
            8'd 97: out = 14'd  169;  // 1/97 ? 0.01030928
            8'd 98: out = 14'd  167;  // 1/98 ? 0.01020408
            8'd 99: out = 14'd  165;  // 1/99 ? 0.01010101
            8'd100: out = 14'd  164;  // 1/100 ? 0.01000000
            8'd101: out = 14'd  162;  // 1/101 ? 0.00990099
            8'd102: out = 14'd  161;  // 1/102 ? 0.00980392
            8'd103: out = 14'd  159;  // 1/103 ? 0.00970874
            8'd104: out = 14'd  158;  // 1/104 ? 0.00961538
            8'd105: out = 14'd  156;  // 1/105 ? 0.00952381
            8'd106: out = 14'd  155;  // 1/106 ? 0.00943396
            8'd107: out = 14'd  153;  // 1/107 ? 0.00934579
            8'd108: out = 14'd  152;  // 1/108 ? 0.00925926
            8'd109: out = 14'd  150;  // 1/109 ? 0.00917431
            8'd110: out = 14'd  149;  // 1/110 ? 0.00909091
            8'd111: out = 14'd  148;  // 1/111 ? 0.00900901
            8'd112: out = 14'd  146;  // 1/112 ? 0.00892857
            8'd113: out = 14'd  145;  // 1/113 ? 0.00884956
            8'd114: out = 14'd  144;  // 1/114 ? 0.00877193
            8'd115: out = 14'd  142;  // 1/115 ? 0.00869565
            8'd116: out = 14'd  141;  // 1/116 ? 0.00862069
            8'd117: out = 14'd  140;  // 1/117 ? 0.00854701
            8'd118: out = 14'd  139;  // 1/118 ? 0.00847458
            8'd119: out = 14'd  138;  // 1/119 ? 0.00840336
            8'd120: out = 14'd  137;  // 1/120 ? 0.00833333
            8'd121: out = 14'd  135;  // 1/121 ? 0.00826446
            8'd122: out = 14'd  134;  // 1/122 ? 0.00819672
            8'd123: out = 14'd  133;  // 1/123 ? 0.00813008
            8'd124: out = 14'd  132;  // 1/124 ? 0.00806452
            8'd125: out = 14'd  131;  // 1/125 ? 0.00800000
            8'd126: out = 14'd  130;  // 1/126 ? 0.00793651
            8'd127: out = 14'd  129;  // 1/127 ? 0.00787402
            8'd128: out = 14'd  128;  // 1/128 ? 0.00781250
            8'd129: out = 14'd  127;  // 1/129 ? 0.00775194
            8'd130: out = 14'd  126;  // 1/130 ? 0.00769231
            8'd131: out = 14'd  125;  // 1/131 ? 0.00763359
            8'd132: out = 14'd  124;  // 1/132 ? 0.00757576
            8'd133: out = 14'd  123;  // 1/133 ? 0.00751880
            8'd134: out = 14'd  122;  // 1/134 ? 0.00746269
            8'd135: out = 14'd  121;  // 1/135 ? 0.00740741
            8'd136: out = 14'd  120;  // 1/136 ? 0.00735294
            8'd137: out = 14'd  120;  // 1/137 ? 0.00729927
            8'd138: out = 14'd  119;  // 1/138 ? 0.00724638
            8'd139: out = 14'd  118;  // 1/139 ? 0.00719424
            8'd140: out = 14'd  117;  // 1/140 ? 0.00714286
            8'd141: out = 14'd  116;  // 1/141 ? 0.00709220
            8'd142: out = 14'd  115;  // 1/142 ? 0.00704225
            8'd143: out = 14'd  115;  // 1/143 ? 0.00699301
            8'd144: out = 14'd  114;  // 1/144 ? 0.00694444
            8'd145: out = 14'd  113;  // 1/145 ? 0.00689655
            8'd146: out = 14'd  112;  // 1/146 ? 0.00684932
            8'd147: out = 14'd  111;  // 1/147 ? 0.00680272
            8'd148: out = 14'd  111;  // 1/148 ? 0.00675676
            8'd149: out = 14'd  110;  // 1/149 ? 0.00671141
            8'd150: out = 14'd  109;  // 1/150 ? 0.00666667
            8'd151: out = 14'd  109;  // 1/151 ? 0.00662252
            8'd152: out = 14'd  108;  // 1/152 ? 0.00657895
            8'd153: out = 14'd  107;  // 1/153 ? 0.00653595
            8'd154: out = 14'd  106;  // 1/154 ? 0.00649351
            8'd155: out = 14'd  106;  // 1/155 ? 0.00645161
            8'd156: out = 14'd  105;  // 1/156 ? 0.00641026
            8'd157: out = 14'd  104;  // 1/157 ? 0.00636943
            8'd158: out = 14'd  104;  // 1/158 ? 0.00632911
            8'd159: out = 14'd  103;  // 1/159 ? 0.00628931
            8'd160: out = 14'd  102;  // 1/160 ? 0.00625000
            8'd161: out = 14'd  102;  // 1/161 ? 0.00621118
            8'd162: out = 14'd  101;  // 1/162 ? 0.00617284
            8'd163: out = 14'd  101;  // 1/163 ? 0.00613497
            8'd164: out = 14'd  100;  // 1/164 ? 0.00609756
            8'd165: out = 14'd   99;  // 1/165 ? 0.00606061
            8'd166: out = 14'd   99;  // 1/166 ? 0.00602410
            8'd167: out = 14'd   98;  // 1/167 ? 0.00598802
            8'd168: out = 14'd   98;  // 1/168 ? 0.00595238
            8'd169: out = 14'd   97;  // 1/169 ? 0.00591716
            8'd170: out = 14'd   96;  // 1/170 ? 0.00588235
            8'd171: out = 14'd   96;  // 1/171 ? 0.00584795
            8'd172: out = 14'd   95;  // 1/172 ? 0.00581395
            8'd173: out = 14'd   95;  // 1/173 ? 0.00578035
            8'd174: out = 14'd   94;  // 1/174 ? 0.00574713
            8'd175: out = 14'd   94;  // 1/175 ? 0.00571429
            8'd176: out = 14'd   93;  // 1/176 ? 0.00568182
            8'd177: out = 14'd   93;  // 1/177 ? 0.00564972
            8'd178: out = 14'd   92;  // 1/178 ? 0.00561798
            8'd179: out = 14'd   92;  // 1/179 ? 0.00558659
            8'd180: out = 14'd   91;  // 1/180 ? 0.00555556
            8'd181: out = 14'd   91;  // 1/181 ? 0.00552486
            8'd182: out = 14'd   90;  // 1/182 ? 0.00549451
            8'd183: out = 14'd   90;  // 1/183 ? 0.00546448
            8'd184: out = 14'd   89;  // 1/184 ? 0.00543478
            8'd185: out = 14'd   89;  // 1/185 ? 0.00540541
            8'd186: out = 14'd   88;  // 1/186 ? 0.00537634
            8'd187: out = 14'd   88;  // 1/187 ? 0.00534759
            8'd188: out = 14'd   87;  // 1/188 ? 0.00531915
            8'd189: out = 14'd   87;  // 1/189 ? 0.00529101
            8'd190: out = 14'd   86;  // 1/190 ? 0.00526316
            8'd191: out = 14'd   86;  // 1/191 ? 0.00523560
            8'd192: out = 14'd   85;  // 1/192 ? 0.00520833
            8'd193: out = 14'd   85;  // 1/193 ? 0.00518135
            8'd194: out = 14'd   84;  // 1/194 ? 0.00515464
            8'd195: out = 14'd   84;  // 1/195 ? 0.00512821
            8'd196: out = 14'd   84;  // 1/196 ? 0.00510204
            8'd197: out = 14'd   83;  // 1/197 ? 0.00507614
            8'd198: out = 14'd   83;  // 1/198 ? 0.00505051
            8'd199: out = 14'd   82;  // 1/199 ? 0.00502513
            8'd200: out = 14'd   82;  // 1/200 ? 0.00500000
            8'd201: out = 14'd   82;  // 1/201 ? 0.00497512
            8'd202: out = 14'd   81;  // 1/202 ? 0.00495050
            8'd203: out = 14'd   81;  // 1/203 ? 0.00492611
            8'd204: out = 14'd   80;  // 1/204 ? 0.00490196
            8'd205: out = 14'd   80;  // 1/205 ? 0.00487805
            8'd206: out = 14'd   80;  // 1/206 ? 0.00485437
            8'd207: out = 14'd   79;  // 1/207 ? 0.00483092
            8'd208: out = 14'd   79;  // 1/208 ? 0.00480769
            8'd209: out = 14'd   78;  // 1/209 ? 0.00478469
            8'd210: out = 14'd   78;  // 1/210 ? 0.00476190
            8'd211: out = 14'd   78;  // 1/211 ? 0.00473934
            8'd212: out = 14'd   77;  // 1/212 ? 0.00471698
            8'd213: out = 14'd   77;  // 1/213 ? 0.00469484
            8'd214: out = 14'd   77;  // 1/214 ? 0.00467290
            8'd215: out = 14'd   76;  // 1/215 ? 0.00465116
            8'd216: out = 14'd   76;  // 1/216 ? 0.00462963
            8'd217: out = 14'd   76;  // 1/217 ? 0.00460829
            8'd218: out = 14'd   75;  // 1/218 ? 0.00458716
            8'd219: out = 14'd   75;  // 1/219 ? 0.00456621
            8'd220: out = 14'd   74;  // 1/220 ? 0.00454545
            8'd221: out = 14'd   74;  // 1/221 ? 0.00452489
            8'd222: out = 14'd   74;  // 1/222 ? 0.00450450
            8'd223: out = 14'd   73;  // 1/223 ? 0.00448430
            8'd224: out = 14'd   73;  // 1/224 ? 0.00446429
            8'd225: out = 14'd   73;  // 1/225 ? 0.00444444
            8'd226: out = 14'd   72;  // 1/226 ? 0.00442478
            8'd227: out = 14'd   72;  // 1/227 ? 0.00440529
            8'd228: out = 14'd   72;  // 1/228 ? 0.00438596
            8'd229: out = 14'd   72;  // 1/229 ? 0.00436681
            8'd230: out = 14'd   71;  // 1/230 ? 0.00434783
            8'd231: out = 14'd   71;  // 1/231 ? 0.00432900
            8'd232: out = 14'd   71;  // 1/232 ? 0.00431034
            8'd233: out = 14'd   70;  // 1/233 ? 0.00429185
            8'd234: out = 14'd   70;  // 1/234 ? 0.00427350
            8'd235: out = 14'd   70;  // 1/235 ? 0.00425532
            8'd236: out = 14'd   69;  // 1/236 ? 0.00423729
            8'd237: out = 14'd   69;  // 1/237 ? 0.00421941
            8'd238: out = 14'd   69;  // 1/238 ? 0.00420168
            8'd239: out = 14'd   69;  // 1/239 ? 0.00418410
            8'd240: out = 14'd   68;  // 1/240 ? 0.00416667
            8'd241: out = 14'd   68;  // 1/241 ? 0.00414938
            8'd242: out = 14'd   68;  // 1/242 ? 0.00413223
            8'd243: out = 14'd   67;  // 1/243 ? 0.00411523
            8'd244: out = 14'd   67;  // 1/244 ? 0.00409836
            8'd245: out = 14'd   67;  // 1/245 ? 0.00408163
            8'd246: out = 14'd   67;  // 1/246 ? 0.00406504
            8'd247: out = 14'd   66;  // 1/247 ? 0.00404858
            8'd248: out = 14'd   66;  // 1/248 ? 0.00403226
            8'd249: out = 14'd   66;  // 1/249 ? 0.00401606
            8'd250: out = 14'd   66;  // 1/250 ? 0.00400000
            8'd251: out = 14'd   65;  // 1/251 ? 0.00398406
            8'd252: out = 14'd   65;  // 1/252 ? 0.00396825
            8'd253: out = 14'd   65;  // 1/253 ? 0.00395257
            8'd254: out = 14'd   65;  // 1/254 ? 0.00393701
            8'd255: out = 14'd   64;  // 1/255 ? 0.00392157
            default: out = 14'd0;  // undefined for 0
        endcase
    end

endmodule
