module Transmission_Reciprocal_LUT (
    input  [9:0] in,      // Q0.10 transmission value (ranges from 0 to 0.65)
    output reg [7:0] out  // Q2.6 reciprocal
);

    always @(*) begin 
        casez (in) 
            10'd   0: out = 8'h40; 
            10'd   1: out = 8'h40;
            10'd   2: out = 8'h40;
            10'd   3: out = 8'h40;
            10'd   4: out = 8'h40;
            10'd   5: out = 8'h40;
            10'd   6: out = 8'h40;
            10'd   7: out = 8'h40;
            10'd   8: out = 8'h41;
            10'd   9: out = 8'h41;
            10'd  10: out = 8'h41;
            10'd  11: out = 8'h41;
            10'd  12: out = 8'h41;
            10'd  13: out = 8'h41;
            10'd  14: out = 8'h41;
            10'd  15: out = 8'h41;
            10'd  16: out = 8'h41;
            10'd  17: out = 8'h41;
            10'd  18: out = 8'h41;
            10'd  19: out = 8'h41;
            10'd  20: out = 8'h41;
            10'd  21: out = 8'h41;
            10'd  22: out = 8'h41;
            10'd  23: out = 8'h41;
            10'd  24: out = 8'h42;
            10'd  25: out = 8'h42;
            10'd  26: out = 8'h42;
            10'd  27: out = 8'h42;
            10'd  28: out = 8'h42;
            10'd  29: out = 8'h42;
            10'd  30: out = 8'h42;
            10'd  31: out = 8'h42;
            10'd  32: out = 8'h42;
            10'd  33: out = 8'h42;
            10'd  34: out = 8'h42;
            10'd  35: out = 8'h42;
            10'd  36: out = 8'h42;
            10'd  37: out = 8'h42;
            10'd  38: out = 8'h42;
            10'd  39: out = 8'h43;
            10'd  40: out = 8'h43;
            10'd  41: out = 8'h43;
            10'd  42: out = 8'h43;
            10'd  43: out = 8'h43;
            10'd  44: out = 8'h43;
            10'd  45: out = 8'h43;
            10'd  46: out = 8'h43;
            10'd  47: out = 8'h43;
            10'd  48: out = 8'h43;
            10'd  49: out = 8'h43;
            10'd  50: out = 8'h43;
            10'd  51: out = 8'h43;
            10'd  52: out = 8'h43;
            10'd  53: out = 8'h43;
            10'd  54: out = 8'h44;
            10'd  55: out = 8'h44;
            10'd  56: out = 8'h44;
            10'd  57: out = 8'h44;
            10'd  58: out = 8'h44;
            10'd  59: out = 8'h44;
            10'd  60: out = 8'h44;
            10'd  61: out = 8'h44;
            10'd  62: out = 8'h44;
            10'd  63: out = 8'h44;
            10'd  64: out = 8'h44;
            10'd  65: out = 8'h44;
            10'd  66: out = 8'h44;
            10'd  67: out = 8'h44;
            10'd  68: out = 8'h45;
            10'd  69: out = 8'h45;
            10'd  70: out = 8'h45;
            10'd  71: out = 8'h45;
            10'd  72: out = 8'h45;
            10'd  73: out = 8'h45;
            10'd  74: out = 8'h45;
            10'd  75: out = 8'h45;
            10'd  76: out = 8'h45;
            10'd  77: out = 8'h45;
            10'd  78: out = 8'h45;
            10'd  79: out = 8'h45;
            10'd  80: out = 8'h45;
            10'd  81: out = 8'h45;
            10'd  82: out = 8'h46;
            10'd  83: out = 8'h46;
            10'd  84: out = 8'h46;
            10'd  85: out = 8'h46;
            10'd  86: out = 8'h46;
            10'd  87: out = 8'h46;
            10'd  88: out = 8'h46;
            10'd  89: out = 8'h46;
            10'd  90: out = 8'h46;
            10'd  91: out = 8'h46;
            10'd  92: out = 8'h46;
            10'd  93: out = 8'h46;
            10'd  94: out = 8'h46;
            10'd  95: out = 8'h47;
            10'd  96: out = 8'h47;
            10'd  97: out = 8'h47;
            10'd  98: out = 8'h47;
            10'd  99: out = 8'h47;
            10'd 100: out = 8'h47;
            10'd 101: out = 8'h47;
            10'd 102: out = 8'h47;
            10'd 103: out = 8'h47;
            10'd 104: out = 8'h47;
            10'd 105: out = 8'h47;
            10'd 106: out = 8'h47;
            10'd 107: out = 8'h47;
            10'd 108: out = 8'h48;
            10'd 109: out = 8'h48;
            10'd 110: out = 8'h48;
            10'd 111: out = 8'h48;
            10'd 112: out = 8'h48;
            10'd 113: out = 8'h48;
            10'd 114: out = 8'h48;
            10'd 115: out = 8'h48;
            10'd 116: out = 8'h48;
            10'd 117: out = 8'h48;
            10'd 118: out = 8'h48;
            10'd 119: out = 8'h48;
            10'd 120: out = 8'h48;
            10'd 121: out = 8'h49;
            10'd 122: out = 8'h49;
            10'd 123: out = 8'h49;
            10'd 124: out = 8'h49;
            10'd 125: out = 8'h49;
            10'd 126: out = 8'h49;
            10'd 127: out = 8'h49;
            10'd 128: out = 8'h49;
            10'd 129: out = 8'h49;
            10'd 130: out = 8'h49;
            10'd 131: out = 8'h49;
            10'd 132: out = 8'h49;
            10'd 133: out = 8'h4A;
            10'd 134: out = 8'h4A;
            10'd 135: out = 8'h4A;
            10'd 136: out = 8'h4A;
            10'd 137: out = 8'h4A;
            10'd 138: out = 8'h4A;
            10'd 139: out = 8'h4A;
            10'd 140: out = 8'h4A;
            10'd 141: out = 8'h4A;
            10'd 142: out = 8'h4A;
            10'd 143: out = 8'h4A;
            10'd 144: out = 8'h4A;
            10'd 145: out = 8'h4B;
            10'd 146: out = 8'h4B;
            10'd 147: out = 8'h4B;
            10'd 148: out = 8'h4B;
            10'd 149: out = 8'h4B;
            10'd 150: out = 8'h4B;
            10'd 151: out = 8'h4B;
            10'd 152: out = 8'h4B;
            10'd 153: out = 8'h4B;
            10'd 154: out = 8'h4B;
            10'd 155: out = 8'h4B;
            10'd 156: out = 8'h4C;
            10'd 157: out = 8'h4C;
            10'd 158: out = 8'h4C;
            10'd 159: out = 8'h4C;
            10'd 160: out = 8'h4C;
            10'd 161: out = 8'h4C;
            10'd 162: out = 8'h4C;
            10'd 163: out = 8'h4C;
            10'd 164: out = 8'h4C;
            10'd 165: out = 8'h4C;
            10'd 166: out = 8'h4C;
            10'd 167: out = 8'h4C;
            10'd 168: out = 8'h4D;
            10'd 169: out = 8'h4D;
            10'd 170: out = 8'h4D;
            10'd 171: out = 8'h4D;
            10'd 172: out = 8'h4D;
            10'd 173: out = 8'h4D;
            10'd 174: out = 8'h4D;
            10'd 175: out = 8'h4D;
            10'd 176: out = 8'h4D;
            10'd 177: out = 8'h4D;
            10'd 178: out = 8'h4D;
            10'd 179: out = 8'h4E;
            10'd 180: out = 8'h4E;
            10'd 181: out = 8'h4E;
            10'd 182: out = 8'h4E;
            10'd 183: out = 8'h4E;
            10'd 184: out = 8'h4E;
            10'd 185: out = 8'h4E;
            10'd 186: out = 8'h4E;
            10'd 187: out = 8'h4E;
            10'd 188: out = 8'h4E;
            10'd 189: out = 8'h4E;
            10'd 190: out = 8'h4F;
            10'd 191: out = 8'h4F;
            10'd 192: out = 8'h4F;
            10'd 193: out = 8'h4F;
            10'd 194: out = 8'h4F;
            10'd 195: out = 8'h4F;
            10'd 196: out = 8'h4F;
            10'd 197: out = 8'h4F;
            10'd 198: out = 8'h4F;
            10'd 199: out = 8'h4F;
            10'd 200: out = 8'h50;
            10'd 201: out = 8'h50;
            10'd 202: out = 8'h50;
            10'd 203: out = 8'h50;
            10'd 204: out = 8'h50;
            10'd 205: out = 8'h50;
            10'd 206: out = 8'h50;
            10'd 207: out = 8'h50;
            10'd 208: out = 8'h50;
            10'd 209: out = 8'h50;
            10'd 210: out = 8'h51;
            10'd 211: out = 8'h51;
            10'd 212: out = 8'h51;
            10'd 213: out = 8'h51;
            10'd 214: out = 8'h51;
            10'd 215: out = 8'h51;
            10'd 216: out = 8'h51;
            10'd 217: out = 8'h51;
            10'd 218: out = 8'h51;
            10'd 219: out = 8'h51;
            10'd 220: out = 8'h52;
            10'd 221: out = 8'h52;
            10'd 222: out = 8'h52;
            10'd 223: out = 8'h52;
            10'd 224: out = 8'h52;
            10'd 225: out = 8'h52;
            10'd 226: out = 8'h52;
            10'd 227: out = 8'h52;
            10'd 228: out = 8'h52;
            10'd 229: out = 8'h52;
            10'd 230: out = 8'h53;
            10'd 231: out = 8'h53;
            10'd 232: out = 8'h53;
            10'd 233: out = 8'h53;
            10'd 234: out = 8'h53;
            10'd 235: out = 8'h53;
            10'd 236: out = 8'h53;
            10'd 237: out = 8'h53;
            10'd 238: out = 8'h53;
            10'd 239: out = 8'h53;
            10'd 240: out = 8'h54;
            10'd 241: out = 8'h54;
            10'd 242: out = 8'h54;
            10'd 243: out = 8'h54;
            10'd 244: out = 8'h54;
            10'd 245: out = 8'h54;
            10'd 246: out = 8'h54;
            10'd 247: out = 8'h54;
            10'd 248: out = 8'h54;
            10'd 249: out = 8'h55;
            10'd 250: out = 8'h55;
            10'd 251: out = 8'h55;
            10'd 252: out = 8'h55;
            10'd 253: out = 8'h55;
            10'd 254: out = 8'h55;
            10'd 255: out = 8'h55;
            10'd 256: out = 8'h55;
            10'd 257: out = 8'h55;
            10'd 258: out = 8'h56;
            10'd 259: out = 8'h56;
            10'd 260: out = 8'h56;
            10'd 261: out = 8'h56;
            10'd 262: out = 8'h56;
            10'd 263: out = 8'h56;
            10'd 264: out = 8'h56;
            10'd 265: out = 8'h56;
            10'd 266: out = 8'h56;
            10'd 267: out = 8'h57;
            10'd 268: out = 8'h57;
            10'd 269: out = 8'h57;
            10'd 270: out = 8'h57;
            10'd 271: out = 8'h57;
            10'd 272: out = 8'h57;
            10'd 273: out = 8'h57;
            10'd 274: out = 8'h57;
            10'd 275: out = 8'h57;
            10'd 276: out = 8'h58;
            10'd 277: out = 8'h58;
            10'd 278: out = 8'h58;
            10'd 279: out = 8'h58;
            10'd 280: out = 8'h58;
            10'd 281: out = 8'h58;
            10'd 282: out = 8'h58;
            10'd 283: out = 8'h58;
            10'd 284: out = 8'h59;
            10'd 285: out = 8'h59;
            10'd 286: out = 8'h59;
            10'd 287: out = 8'h59;
            10'd 288: out = 8'h59;
            10'd 289: out = 8'h59;
            10'd 290: out = 8'h59;
            10'd 291: out = 8'h59;
            10'd 292: out = 8'h5A;
            10'd 293: out = 8'h5A;
            10'd 294: out = 8'h5A;
            10'd 295: out = 8'h5A;
            10'd 296: out = 8'h5A;
            10'd 297: out = 8'h5A;
            10'd 298: out = 8'h5A;
            10'd 299: out = 8'h5A;
            10'd 300: out = 8'h5B;
            10'd 301: out = 8'h5B;
            10'd 302: out = 8'h5B;
            10'd 303: out = 8'h5B;
            10'd 304: out = 8'h5B;
            10'd 305: out = 8'h5B;
            10'd 306: out = 8'h5B;
            10'd 307: out = 8'h5B;
            10'd 308: out = 8'h5C;
            10'd 309: out = 8'h5C;
            10'd 310: out = 8'h5C;
            10'd 311: out = 8'h5C;
            10'd 312: out = 8'h5C;
            10'd 313: out = 8'h5C;
            10'd 314: out = 8'h5C;
            10'd 315: out = 8'h5C;
            10'd 316: out = 8'h5D;
            10'd 317: out = 8'h5D;
            10'd 318: out = 8'h5D;
            10'd 319: out = 8'h5D;
            10'd 320: out = 8'h5D;
            10'd 321: out = 8'h5D;
            10'd 322: out = 8'h5D;
            10'd 323: out = 8'h5D;
            10'd 324: out = 8'h5E;
            10'd 325: out = 8'h5E;
            10'd 326: out = 8'h5E;
            10'd 327: out = 8'h5E;
            10'd 328: out = 8'h5E;
            10'd 329: out = 8'h5E;
            10'd 330: out = 8'h5E;
            10'd 331: out = 8'h5F;
            10'd 332: out = 8'h5F;
            10'd 333: out = 8'h5F;
            10'd 334: out = 8'h5F;
            10'd 335: out = 8'h5F;
            10'd 336: out = 8'h5F;
            10'd 337: out = 8'h5F;
            10'd 338: out = 8'h60;
            10'd 339: out = 8'h60;
            10'd 340: out = 8'h60;
            10'd 341: out = 8'h60;
            10'd 342: out = 8'h60;
            10'd 343: out = 8'h60;
            10'd 344: out = 8'h60;
            10'd 345: out = 8'h61;
            10'd 346: out = 8'h61;
            10'd 347: out = 8'h61;
            10'd 348: out = 8'h61;
            10'd 349: out = 8'h61;
            10'd 350: out = 8'h61;
            10'd 351: out = 8'h61;
            10'd 352: out = 8'h62;
            10'd 353: out = 8'h62;
            10'd 354: out = 8'h62;
            10'd 355: out = 8'h62;
            10'd 356: out = 8'h62;
            10'd 357: out = 8'h62;
            10'd 358: out = 8'h62;
            10'd 359: out = 8'h63;
            10'd 360: out = 8'h63;
            10'd 361: out = 8'h63;
            10'd 362: out = 8'h63;
            10'd 363: out = 8'h63;
            10'd 364: out = 8'h63;
            10'd 365: out = 8'h63;
            10'd 366: out = 8'h64;
            10'd 367: out = 8'h64;
            10'd 368: out = 8'h64;
            10'd 369: out = 8'h64;
            10'd 370: out = 8'h64;
            10'd 371: out = 8'h64;
            10'd 372: out = 8'h65;
            10'd 373: out = 8'h65;
            10'd 374: out = 8'h65;
            10'd 375: out = 8'h65;
            10'd 376: out = 8'h65;
            10'd 377: out = 8'h65;
            10'd 378: out = 8'h65;
            10'd 379: out = 8'h66;
            10'd 380: out = 8'h66;
            10'd 381: out = 8'h66;
            10'd 382: out = 8'h66;
            10'd 383: out = 8'h66;
            10'd 384: out = 8'h66;
            10'd 385: out = 8'h67;
            10'd 386: out = 8'h67;
            10'd 387: out = 8'h67;
            10'd 388: out = 8'h67;
            10'd 389: out = 8'h67;
            10'd 390: out = 8'h67;
            10'd 391: out = 8'h68;
            10'd 392: out = 8'h68;
            10'd 393: out = 8'h68;
            10'd 394: out = 8'h68;
            10'd 395: out = 8'h68;
            10'd 396: out = 8'h68;
            10'd 397: out = 8'h69;
            10'd 398: out = 8'h69;
            10'd 399: out = 8'h69;
            10'd 400: out = 8'h69;
            10'd 401: out = 8'h69;
            10'd 402: out = 8'h69;
            10'd 403: out = 8'h6A;
            10'd 404: out = 8'h6A;
            10'd 405: out = 8'h6A;
            10'd 406: out = 8'h6A;
            10'd 407: out = 8'h6A;
            10'd 408: out = 8'h6A;
            10'd 409: out = 8'h6B;
            10'd 410: out = 8'h6B;
            10'd 411: out = 8'h6B;
            10'd 412: out = 8'h6B;
            10'd 413: out = 8'h6B;
            10'd 414: out = 8'h6B;
            10'd 415: out = 8'h6C;
            10'd 416: out = 8'h6C;
            10'd 417: out = 8'h6C;
            10'd 418: out = 8'h6C;
            10'd 419: out = 8'h6C;
            10'd 420: out = 8'h6D;
            10'd 421: out = 8'h6D;
            10'd 422: out = 8'h6D;
            10'd 423: out = 8'h6D;
            10'd 424: out = 8'h6D;
            10'd 425: out = 8'h6D;
            10'd 426: out = 8'h6E;
            10'd 427: out = 8'h6E;
            10'd 428: out = 8'h6E;
            10'd 429: out = 8'h6E;
            10'd 430: out = 8'h6E;
            10'd 431: out = 8'h6F;
            10'd 432: out = 8'h6F;
            10'd 433: out = 8'h6F;
            10'd 434: out = 8'h6F;
            10'd 435: out = 8'h6F;
            10'd 436: out = 8'h6F;
            10'd 437: out = 8'h70;
            10'd 438: out = 8'h70;
            10'd 439: out = 8'h70;
            10'd 440: out = 8'h70;
            10'd 441: out = 8'h70;
            10'd 442: out = 8'h71;
            10'd 443: out = 8'h71;
            10'd 444: out = 8'h71;
            10'd 445: out = 8'h71;
            10'd 446: out = 8'h71;
            10'd 447: out = 8'h72;
            10'd 448: out = 8'h72;
            10'd 449: out = 8'h72;
            10'd 450: out = 8'h72;
            10'd 451: out = 8'h72;
            10'd 452: out = 8'h73;
            10'd 453: out = 8'h73;
            10'd 454: out = 8'h73;
            10'd 455: out = 8'h73;
            10'd 456: out = 8'h73;
            10'd 457: out = 8'h74;
            10'd 458: out = 8'h74;
            10'd 459: out = 8'h74;
            10'd 460: out = 8'h74;
            10'd 461: out = 8'h74;
            10'd 462: out = 8'h75;
            10'd 463: out = 8'h75;
            10'd 464: out = 8'h75;
            10'd 465: out = 8'h75;
            10'd 466: out = 8'h75;
            10'd 467: out = 8'h76;
            10'd 468: out = 8'h76;
            10'd 469: out = 8'h76;
            10'd 470: out = 8'h76;
            10'd 471: out = 8'h77;
            10'd 472: out = 8'h77;
            10'd 473: out = 8'h77;
            10'd 474: out = 8'h77;
            10'd 475: out = 8'h77;
            10'd 476: out = 8'h78;
            10'd 477: out = 8'h78;
            10'd 478: out = 8'h78;
            10'd 479: out = 8'h78;
            10'd 480: out = 8'h78;
            10'd 481: out = 8'h79;
            10'd 482: out = 8'h79;
            10'd 483: out = 8'h79;
            10'd 484: out = 8'h79;
            10'd 485: out = 8'h7A;
            10'd 486: out = 8'h7A;
            10'd 487: out = 8'h7A;
            10'd 488: out = 8'h7A;
            10'd 489: out = 8'h7A;
            10'd 490: out = 8'h7B;
            10'd 491: out = 8'h7B;
            10'd 492: out = 8'h7B;
            10'd 493: out = 8'h7B;
            10'd 494: out = 8'h7C;
            10'd 495: out = 8'h7C;
            10'd 496: out = 8'h7C;
            10'd 497: out = 8'h7C;
            10'd 498: out = 8'h7D;
            10'd 499: out = 8'h7D;
            10'd 500: out = 8'h7D;
            10'd 501: out = 8'h7D;
            10'd 502: out = 8'h7E;
            10'd 503: out = 8'h7E;
            10'd 504: out = 8'h7E;
            10'd 505: out = 8'h7E;
            10'd 506: out = 8'h7F;
            10'd 507: out = 8'h7F;
            10'd 508: out = 8'h7F;
            10'd 509: out = 8'h7F;
            10'd 510: out = 8'h80;
            10'd 511: out = 8'h80;
            10'd 512: out = 8'h80;
            10'd 513: out = 8'h80;
            10'd 514: out = 8'h81;
            10'd 515: out = 8'h81;
            10'd 516: out = 8'h81;
            10'd 517: out = 8'h81;
            10'd 518: out = 8'h82;
            10'd 519: out = 8'h82;
            10'd 520: out = 8'h82;
            10'd 521: out = 8'h82;
            10'd 522: out = 8'h83;
            10'd 523: out = 8'h83;
            10'd 524: out = 8'h83;
            10'd 525: out = 8'h83;
            10'd 526: out = 8'h84;
            10'd 527: out = 8'h84;
            10'd 528: out = 8'h84;
            10'd 529: out = 8'h84;
            10'd 530: out = 8'h85;
            10'd 531: out = 8'h85;
            10'd 532: out = 8'h85;
            10'd 533: out = 8'h85;
            10'd 534: out = 8'h86;
            10'd 535: out = 8'h86;
            10'd 536: out = 8'h86;
            10'd 537: out = 8'h87;
            10'd 538: out = 8'h87;
            10'd 539: out = 8'h87;
            10'd 540: out = 8'h87;
            10'd 541: out = 8'h88;
            10'd 542: out = 8'h88;
            10'd 543: out = 8'h88;
            10'd 544: out = 8'h89;
            10'd 545: out = 8'h89;
            10'd 546: out = 8'h89;
            10'd 547: out = 8'h89;
            10'd 548: out = 8'h8A;
            10'd 549: out = 8'h8A;
            10'd 550: out = 8'h8A;
            10'd 551: out = 8'h8B;
            10'd 552: out = 8'h8B;
            10'd 553: out = 8'h8B;
            10'd 554: out = 8'h8B;
            10'd 555: out = 8'h8C;
            10'd 556: out = 8'h8C;
            10'd 557: out = 8'h8C;
            10'd 558: out = 8'h8D;
            10'd 559: out = 8'h8D;
            10'd 560: out = 8'h8D;
            10'd 561: out = 8'h8E;
            10'd 562: out = 8'h8E;
            10'd 563: out = 8'h8E;
            10'd 564: out = 8'h8E;
            10'd 565: out = 8'h8F;
            10'd 566: out = 8'h8F;
            10'd 567: out = 8'h8F;
            10'd 568: out = 8'h90;
            10'd 569: out = 8'h90;
            10'd 570: out = 8'h90;
            10'd 571: out = 8'h91;
            10'd 572: out = 8'h91;
            10'd 573: out = 8'h91;
            10'd 574: out = 8'h92;
            10'd 575: out = 8'h92;
            10'd 576: out = 8'h92;
            10'd 577: out = 8'h93;
            10'd 578: out = 8'h93;
            10'd 579: out = 8'h93;
            10'd 580: out = 8'h94;
            10'd 581: out = 8'h94;
            10'd 582: out = 8'h94;
            10'd 583: out = 8'h95;
            10'd 584: out = 8'h95;
            10'd 585: out = 8'h95;
            10'd 586: out = 8'h96;
            10'd 587: out = 8'h96;
            10'd 588: out = 8'h96;
            10'd 589: out = 8'h97;
            10'd 590: out = 8'h97;
            10'd 591: out = 8'h97;
            10'd 592: out = 8'h98;
            10'd 593: out = 8'h98;
            10'd 594: out = 8'h98;
            10'd 595: out = 8'h99;
            10'd 596: out = 8'h99;
            10'd 597: out = 8'h99;
            10'd 598: out = 8'h9A;
            10'd 599: out = 8'h9A;
            10'd 600: out = 8'h9B;
            10'd 601: out = 8'h9B;
            10'd 602: out = 8'h9B;
            10'd 603: out = 8'h9C;
            10'd 604: out = 8'h9C;
            10'd 605: out = 8'h9C;
            10'd 606: out = 8'h9D;
            10'd 607: out = 8'h9D;
            10'd 608: out = 8'h9E;
            10'd 609: out = 8'h9E;
            10'd 610: out = 8'h9E;
            10'd 611: out = 8'h9F;
            10'd 612: out = 8'h9F;
            10'd 613: out = 8'h9F;
            10'd 614: out = 8'hA0;
            10'd 615: out = 8'hA0;
            10'd 616: out = 8'hA1;
            10'd 617: out = 8'hA1;
            10'd 618: out = 8'hA1;
            10'd 619: out = 8'hA2;
            10'd 620: out = 8'hA2;
            10'd 621: out = 8'hA3;
            10'd 622: out = 8'hA3;
            10'd 623: out = 8'hA3;
            10'd 624: out = 8'hA4;
            10'd 625: out = 8'hA4;
            10'd 626: out = 8'hA5;
            10'd 627: out = 8'hA5;
            10'd 628: out = 8'hA5;
            10'd 629: out = 8'hA6;
            10'd 630: out = 8'hA6;
            10'd 631: out = 8'hA7;
            10'd 632: out = 8'hA7;
            10'd 633: out = 8'hA8;
            10'd 634: out = 8'hA8;
            10'd 635: out = 8'hA8;
            10'd 636: out = 8'hA9;
            10'd 637: out = 8'hA9;
            10'd 638: out = 8'hAA;
            10'd 639: out = 8'hAA;
            10'd 640: out = 8'hAB;
            10'd 641: out = 8'hAB;
            10'd 642: out = 8'hAC;
            10'd 643: out = 8'hAC;
            10'd 644: out = 8'hAC;
            10'd 645: out = 8'hAD;
            10'd 646: out = 8'hAD;
            10'd 647: out = 8'hAE;
            10'd 648: out = 8'hAE;
            10'd 649: out = 8'hAF;
            10'd 650: out = 8'hAF;
            10'd 651: out = 8'hB0;
            10'd 652: out = 8'hB0;
            10'd 653: out = 8'hB1;
            10'd 654: out = 8'hB1;
            10'd 655: out = 8'hB2;
            10'd 656: out = 8'hB2;
            10'd 657: out = 8'hB3;
            10'd 658: out = 8'hB3;
            10'd 659: out = 8'hB4;
            10'd 660: out = 8'hB4;
            10'd 661: out = 8'hB5;
            10'd 662: out = 8'hB5;
            10'd 663: out = 8'hB6;
            10'd 664: out = 8'hB6;
            10'd 665: out = 8'hB7;
            10'd 666: out = 8'hB7;
            default:  out = 8'hB8;
        endcase
    end
endmodule
