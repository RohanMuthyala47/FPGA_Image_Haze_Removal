// LUT for x^0.3 in Q3.7 format
module LUT_03 (
    input      [7:0] in, // Q8.0 input
    output reg [9:0] out // Q3.7 output
);

    always @(*) begin
        casez (in)
            8'd0  : out = 10'd0;  // 0^0.30 ~= 0.000000
            8'd1  : out = 10'd128;  // 1^0.30 ~= 1.000000
            8'd2  : out = 10'd158;  // 2^0.30 ~= 1.231144
            8'd3  : out = 10'd178;  // 3^0.30 ~= 1.390389
            8'd4  : out = 10'd194;  // 4^0.30 ~= 1.515717
            8'd5  : out = 10'd207;  // 5^0.30 ~= 1.620657
            8'd6  : out = 10'd219;  // 6^0.30 ~= 1.711770
            8'd7  : out = 10'd229;  // 7^0.30 ~= 1.792790
            8'd8  : out = 10'd239;  // 8^0.30 ~= 1.866066
            8'd9  : out = 10'd247;  // 9^0.30 ~= 1.933182
            8'd10 : out = 10'd255;  // 10^0.30 ~= 1.995262
            8'd11 : out = 10'd263;  // 11^0.30 ~= 2.053136
            8'd12 : out = 10'd270;  // 12^0.30 ~= 2.107436
            8'd13 : out = 10'd276;  // 13^0.30 ~= 2.158654
            8'd14 : out = 10'd283;  // 14^0.30 ~= 2.207183
            8'd15 : out = 10'd288;  // 15^0.30 ~= 2.253343
            8'd16 : out = 10'd294;  // 16^0.30 ~= 2.297397
            8'd17 : out = 10'd299;  // 17^0.30 ~= 2.339563
            8'd18 : out = 10'd305;  // 18^0.30 ~= 2.380026
            8'd19 : out = 10'd310;  // 19^0.30 ~= 2.418945
            8'd20 : out = 10'd314;  // 20^0.30 ~= 2.456456
            8'd21 : out = 10'd319;  // 21^0.30 ~= 2.492676
            8'd22 : out = 10'd324;  // 22^0.30 ~= 2.527707
            8'd23 : out = 10'd328;  // 23^0.30 ~= 2.561642
            8'd24 : out = 10'd332;  // 24^0.30 ~= 2.594558
            8'd25 : out = 10'd336;  // 25^0.30 ~= 2.626528
            8'd26 : out = 10'd340;  // 26^0.30 ~= 2.657615
            8'd27 : out = 10'd344;  // 27^0.30 ~= 2.687875
            8'd28 : out = 10'd348;  // 28^0.30 ~= 2.717361
            8'd29 : out = 10'd352;  // 29^0.30 ~= 2.746119
            8'd30 : out = 10'd355;  // 30^0.30 ~= 2.774191
            8'd31 : out = 10'd359;  // 31^0.30 ~= 2.801615
            8'd32 : out = 10'd362;  // 32^0.30 ~= 2.828427
            8'd33 : out = 10'd365;  // 33^0.30 ~= 2.854659
            8'd34 : out = 10'd369;  // 34^0.30 ~= 2.880339
            8'd35 : out = 10'd372;  // 35^0.30 ~= 2.905497
            8'd36 : out = 10'd375;  // 36^0.30 ~= 2.930156
            8'd37 : out = 10'd378;  // 37^0.30 ~= 2.954340
            8'd38 : out = 10'd381;  // 38^0.30 ~= 2.978071
            8'd39 : out = 10'd384;  // 39^0.30 ~= 3.001369
            8'd40 : out = 10'd387;  // 40^0.30 ~= 3.024252
            8'd41 : out = 10'd390;  // 41^0.30 ~= 3.046738
            8'd42 : out = 10'd393;  // 42^0.30 ~= 3.068844
            8'd43 : out = 10'd396;  // 43^0.30 ~= 3.090584
            8'd44 : out = 10'd398;  // 44^0.30 ~= 3.111973
            8'd45 : out = 10'd401;  // 45^0.30 ~= 3.133024
            8'd46 : out = 10'd404;  // 46^0.30 ~= 3.153751
            8'd47 : out = 10'd406;  // 47^0.30 ~= 3.174164
            8'd48 : out = 10'd409;  // 48^0.30 ~= 3.194276
            8'd49 : out = 10'd411;  // 49^0.30 ~= 3.214096
            8'd50 : out = 10'd414;  // 50^0.30 ~= 3.233635
            8'd51 : out = 10'd416;  // 51^0.30 ~= 3.252903
            8'd52 : out = 10'd419;  // 52^0.30 ~= 3.271907
            8'd53 : out = 10'd421;  // 53^0.30 ~= 3.290658
            8'd54 : out = 10'd424;  // 54^0.30 ~= 3.309163
            8'd55 : out = 10'd426;  // 55^0.30 ~= 3.327429
            8'd56 : out = 10'd428;  // 56^0.30 ~= 3.345464
            8'd57 : out = 10'd430;  // 57^0.30 ~= 3.363276
            8'd58 : out = 10'd433;  // 58^0.30 ~= 3.380869
            8'd59 : out = 10'd435;  // 59^0.30 ~= 3.398252
            8'd60 : out = 10'd437;  // 60^0.30 ~= 3.415430
            8'd61 : out = 10'd439;  // 61^0.30 ~= 3.432408
            8'd62 : out = 10'd441;  // 62^0.30 ~= 3.449193
            8'd63 : out = 10'd444;  // 63^0.30 ~= 3.465789
            8'd64 : out = 10'd446;  // 64^0.30 ~= 3.482202
            8'd65 : out = 10'd448;  // 65^0.30 ~= 3.498437
            8'd66 : out = 10'd450;  // 66^0.30 ~= 3.514497
            8'd67 : out = 10'd452;  // 67^0.30 ~= 3.530388
            8'd68 : out = 10'd454;  // 68^0.30 ~= 3.546114
            8'd69 : out = 10'd456;  // 69^0.30 ~= 3.561679
            8'd70 : out = 10'd458;  // 70^0.30 ~= 3.577086
            8'd71 : out = 10'd460;  // 71^0.30 ~= 3.592341
            8'd72 : out = 10'd462;  // 72^0.30 ~= 3.607445
            8'd73 : out = 10'd464;  // 73^0.30 ~= 3.622404
            8'd74 : out = 10'd466;  // 74^0.30 ~= 3.637220
            8'd75 : out = 10'd467;  // 75^0.30 ~= 3.651896
            8'd76 : out = 10'd469;  // 76^0.30 ~= 3.666436
            8'd77 : out = 10'd471;  // 77^0.30 ~= 3.680842
            8'd78 : out = 10'd473;  // 78^0.30 ~= 3.695119
            8'd79 : out = 10'd475;  // 79^0.30 ~= 3.709267
            8'd80 : out = 10'd477;  // 80^0.30 ~= 3.723291
            8'd81 : out = 10'd478;  // 81^0.30 ~= 3.737193
            8'd82 : out = 10'd480;  // 82^0.30 ~= 3.750975
            8'd83 : out = 10'd482;  // 83^0.30 ~= 3.764640
            8'd84 : out = 10'd484;  // 84^0.30 ~= 3.778190
            8'd85 : out = 10'd485;  // 85^0.30 ~= 3.791628
            8'd86 : out = 10'd487;  // 86^0.30 ~= 3.804955
            8'd87 : out = 10'd489;  // 87^0.30 ~= 3.818175
            8'd88 : out = 10'd490;  // 88^0.30 ~= 3.831288
            8'd89 : out = 10'd492;  // 89^0.30 ~= 3.844298
            8'd90 : out = 10'd494;  // 90^0.30 ~= 3.857205
            8'd91 : out = 10'd495;  // 91^0.30 ~= 3.870013
            8'd92 : out = 10'd497;  // 92^0.30 ~= 3.882722
            8'd93 : out = 10'd499;  // 93^0.30 ~= 3.895336
            8'd94 : out = 10'd500;  // 94^0.30 ~= 3.907854
            8'd95 : out = 10'd502;  // 95^0.30 ~= 3.920280
            8'd96 : out = 10'd503;  // 96^0.30 ~= 3.932614
            8'd97 : out = 10'd505;  // 97^0.30 ~= 3.944859
            8'd98 : out = 10'd506;  // 98^0.30 ~= 3.957016
            8'd99 : out = 10'd508;  // 99^0.30 ~= 3.969086
            8'd100: out = 10'd510;  // 100^0.30 ~= 3.981072
            8'd101: out = 10'd511;  // 101^0.30 ~= 3.992973
            8'd102: out = 10'd513;  // 102^0.30 ~= 4.004793
            8'd103: out = 10'd514;  // 103^0.30 ~= 4.016531
            8'd104: out = 10'd516;  // 104^0.30 ~= 4.028191
            8'd105: out = 10'd517;  // 105^0.30 ~= 4.039771
            8'd106: out = 10'd519;  // 106^0.30 ~= 4.051275
            8'd107: out = 10'd520;  // 107^0.30 ~= 4.062704
            8'd108: out = 10'd521;  // 108^0.30 ~= 4.074057
            8'd109: out = 10'd523;  // 109^0.30 ~= 4.085338
            8'd110: out = 10'd524;  // 110^0.30 ~= 4.096546
            8'd111: out = 10'd526;  // 111^0.30 ~= 4.107683
            8'd112: out = 10'd527;  // 112^0.30 ~= 4.118750
            8'd113: out = 10'd529;  // 113^0.30 ~= 4.129748
            8'd114: out = 10'd530;  // 114^0.30 ~= 4.140678
            8'd115: out = 10'd531;  // 115^0.30 ~= 4.151541
            8'd116: out = 10'd533;  // 116^0.30 ~= 4.162339
            8'd117: out = 10'd534;  // 117^0.30 ~= 4.173071
            8'd118: out = 10'd536;  // 118^0.30 ~= 4.183739
            8'd119: out = 10'd537;  // 119^0.30 ~= 4.194344
            8'd120: out = 10'd538;  // 120^0.30 ~= 4.204887
            8'd121: out = 10'd540;  // 121^0.30 ~= 4.215369
            8'd122: out = 10'd541;  // 122^0.30 ~= 4.225790
            8'd123: out = 10'd542;  // 123^0.30 ~= 4.236152
            8'd124: out = 10'd544;  // 124^0.30 ~= 4.246455
            8'd125: out = 10'd545;  // 125^0.30 ~= 4.256700
            8'd126: out = 10'd546;  // 126^0.30 ~= 4.266887
            8'd127: out = 10'd547;  // 127^0.30 ~= 4.277018
            8'd128: out = 10'd549;  // 128^0.30 ~= 4.287094
            8'd129: out = 10'd550;  // 129^0.30 ~= 4.297114
            8'd130: out = 10'd551;  // 130^0.30 ~= 4.307081
            8'd131: out = 10'd553;  // 131^0.30 ~= 4.316993
            8'd132: out = 10'd554;  // 132^0.30 ~= 4.326853
            8'd133: out = 10'd555;  // 133^0.30 ~= 4.336661
            8'd134: out = 10'd556;  // 134^0.30 ~= 4.346417
            8'd135: out = 10'd558;  // 135^0.30 ~= 4.356123
            8'd136: out = 10'd559;  // 136^0.30 ~= 4.365778
            8'd137: out = 10'd560;  // 137^0.30 ~= 4.375384
            8'd138: out = 10'd561;  // 138^0.30 ~= 4.384941
            8'd139: out = 10'd562;  // 139^0.30 ~= 4.394449
            8'd140: out = 10'd564;  // 140^0.30 ~= 4.403910
            8'd141: out = 10'd565;  // 141^0.30 ~= 4.413323
            8'd142: out = 10'd566;  // 142^0.30 ~= 4.422690
            8'd143: out = 10'd567;  // 143^0.30 ~= 4.432011
            8'd144: out = 10'd568;  // 144^0.30 ~= 4.441286
            8'd145: out = 10'd570;  // 145^0.30 ~= 4.450516
            8'd146: out = 10'd571;  // 146^0.30 ~= 4.459702
            8'd147: out = 10'd572;  // 147^0.30 ~= 4.468844
            8'd148: out = 10'd573;  // 148^0.30 ~= 4.477943
            8'd149: out = 10'd574;  // 149^0.30 ~= 4.486998
            8'd150: out = 10'd575;  // 150^0.30 ~= 4.496011
            8'd151: out = 10'd577;  // 151^0.30 ~= 4.504982
            8'd152: out = 10'd578;  // 152^0.30 ~= 4.513912
            8'd153: out = 10'd579;  // 153^0.30 ~= 4.522800
            8'd154: out = 10'd580;  // 154^0.30 ~= 4.531649
            8'd155: out = 10'd581;  // 155^0.30 ~= 4.540456
            8'd156: out = 10'd582;  // 156^0.30 ~= 4.549225
            8'd157: out = 10'd583;  // 157^0.30 ~= 4.557954
            8'd158: out = 10'd585;  // 158^0.30 ~= 4.566644
            8'd159: out = 10'd586;  // 159^0.30 ~= 4.575295
            8'd160: out = 10'd587;  // 160^0.30 ~= 4.583909
            8'd161: out = 10'd588;  // 161^0.30 ~= 4.592485
            8'd162: out = 10'd589;  // 162^0.30 ~= 4.601024
            8'd163: out = 10'd590;  // 163^0.30 ~= 4.609526
            8'd164: out = 10'd591;  // 164^0.30 ~= 4.617992
            8'd165: out = 10'd592;  // 165^0.30 ~= 4.626421
            8'd166: out = 10'd593;  // 166^0.30 ~= 4.634815
            8'd167: out = 10'd594;  // 167^0.30 ~= 4.643174
            8'd168: out = 10'd595;  // 168^0.30 ~= 4.651497
            8'd169: out = 10'd596;  // 169^0.30 ~= 4.659786
            8'd170: out = 10'd598;  // 170^0.30 ~= 4.668041
            8'd171: out = 10'd599;  // 171^0.30 ~= 4.676262
            8'd172: out = 10'd600;  // 172^0.30 ~= 4.684449
            8'd173: out = 10'd601;  // 173^0.30 ~= 4.692603
            8'd174: out = 10'd602;  // 174^0.30 ~= 4.700724
            8'd175: out = 10'd603;  // 175^0.30 ~= 4.708813
            8'd176: out = 10'd604;  // 176^0.30 ~= 4.716869
            8'd177: out = 10'd605;  // 177^0.30 ~= 4.724893
            8'd178: out = 10'd606;  // 178^0.30 ~= 4.732886
            8'd179: out = 10'd607;  // 179^0.30 ~= 4.740847
            8'd180: out = 10'd608;  // 180^0.30 ~= 4.748777
            8'd181: out = 10'd609;  // 181^0.30 ~= 4.756676
            8'd182: out = 10'd610;  // 182^0.30 ~= 4.764545
            8'd183: out = 10'd611;  // 183^0.30 ~= 4.772383
            8'd184: out = 10'd612;  // 184^0.30 ~= 4.780192
            8'd185: out = 10'd613;  // 185^0.30 ~= 4.787971
            8'd186: out = 10'd614;  // 186^0.30 ~= 4.795721
            8'd187: out = 10'd615;  // 187^0.30 ~= 4.803441
            8'd188: out = 10'd616;  // 188^0.30 ~= 4.811133
            8'd189: out = 10'd617;  // 189^0.30 ~= 4.818796
            8'd190: out = 10'd618;  // 190^0.30 ~= 4.826431
            8'd191: out = 10'd619;  // 191^0.30 ~= 4.834037
            8'd192: out = 10'd620;  // 192^0.30 ~= 4.841616
            8'd193: out = 10'd621;  // 193^0.30 ~= 4.849168
            8'd194: out = 10'd622;  // 194^0.30 ~= 4.856692
            8'd195: out = 10'd623;  // 195^0.30 ~= 4.864188
            8'd196: out = 10'd624;  // 196^0.30 ~= 4.871658
            8'd197: out = 10'd625;  // 197^0.30 ~= 4.879102
            8'd198: out = 10'd625;  // 198^0.30 ~= 4.886519
            8'd199: out = 10'd626;  // 199^0.30 ~= 4.893909
            8'd200: out = 10'd627;  // 200^0.30 ~= 4.901274
            8'd201: out = 10'd628;  // 201^0.30 ~= 4.908613
            8'd202: out = 10'd629;  // 202^0.30 ~= 4.915927
            8'd203: out = 10'd630;  // 203^0.30 ~= 4.923215
            8'd204: out = 10'd631;  // 204^0.30 ~= 4.930478
            8'd205: out = 10'd632;  // 205^0.30 ~= 4.937717
            8'd206: out = 10'd633;  // 206^0.30 ~= 4.944930
            8'd207: out = 10'd634;  // 207^0.30 ~= 4.952119
            8'd208: out = 10'd635;  // 208^0.30 ~= 4.959284
            8'd209: out = 10'd636;  // 209^0.30 ~= 4.966425
            8'd210: out = 10'd637;  // 210^0.30 ~= 4.973542
            8'd211: out = 10'd638;  // 211^0.30 ~= 4.980635
            8'd212: out = 10'd638;  // 212^0.30 ~= 4.987705
            8'd213: out = 10'd639;  // 213^0.30 ~= 4.994751
            8'd214: out = 10'd640;  // 214^0.30 ~= 5.001775
            8'd215: out = 10'd641;  // 215^0.30 ~= 5.008775
            8'd216: out = 10'd642;  // 216^0.30 ~= 5.015753
            8'd217: out = 10'd643;  // 217^0.30 ~= 5.022708
            8'd218: out = 10'd644;  // 218^0.30 ~= 5.029641
            8'd219: out = 10'd645;  // 219^0.30 ~= 5.036551
            8'd220: out = 10'd646;  // 220^0.30 ~= 5.043439
            8'd221: out = 10'd646;  // 221^0.30 ~= 5.050306
            8'd222: out = 10'd647;  // 222^0.30 ~= 5.057151
            8'd223: out = 10'd648;  // 223^0.30 ~= 5.063974
            8'd224: out = 10'd649;  // 224^0.30 ~= 5.070776
            8'd225: out = 10'd650;  // 225^0.30 ~= 5.077556
            8'd226: out = 10'd651;  // 226^0.30 ~= 5.084316
            8'd227: out = 10'd652;  // 227^0.30 ~= 5.091055
            8'd228: out = 10'd653;  // 228^0.30 ~= 5.097773
            8'd229: out = 10'd653;  // 229^0.30 ~= 5.104470
            8'd230: out = 10'd654;  // 230^0.30 ~= 5.111147
            8'd231: out = 10'd655;  // 231^0.30 ~= 5.117803
            8'd232: out = 10'd656;  // 232^0.30 ~= 5.124440
            8'd233: out = 10'd657;  // 233^0.30 ~= 5.131056
            8'd234: out = 10'd658;  // 234^0.30 ~= 5.137653
            8'd235: out = 10'd658;  // 235^0.30 ~= 5.144230
            8'd236: out = 10'd659;  // 236^0.30 ~= 5.150787
            8'd237: out = 10'd660;  // 237^0.30 ~= 5.157325
            8'd238: out = 10'd661;  // 238^0.30 ~= 5.163844
            8'd239: out = 10'd662;  // 239^0.30 ~= 5.170343
            8'd240: out = 10'd663;  // 240^0.30 ~= 5.176824
            8'd241: out = 10'd663;  // 241^0.30 ~= 5.183285
            8'd242: out = 10'd664;  // 242^0.30 ~= 5.189728
            8'd243: out = 10'd665;  // 243^0.30 ~= 5.196152
            8'd244: out = 10'd666;  // 244^0.30 ~= 5.202558
            8'd245: out = 10'd667;  // 245^0.30 ~= 5.208946
            8'd246: out = 10'd668;  // 246^0.30 ~= 5.215315
            8'd247: out = 10'd668;  // 247^0.30 ~= 5.221666
            8'd248: out = 10'd669;  // 248^0.30 ~= 5.227999
            8'd249: out = 10'd670;  // 249^0.30 ~= 5.234314
            8'd250: out = 10'd671;  // 250^0.30 ~= 5.240612
            8'd251: out = 10'd672;  // 251^0.30 ~= 5.246892
            8'd252: out = 10'd672;  // 252^0.30 ~= 5.253154
            8'd253: out = 10'd673;  // 253^0.30 ~= 5.259399
            8'd254: out = 10'd674;  // 254^0.30 ~= 5.265627
            8'd255: out = 10'd675;  // 255^0.30 ~= 5.271838
            default: out = 10'd0;
        endcase
    end
endmodule


// LUT for x^0.7 in Q6.4 format
module LUT_07 (
    input      [7:0] in, // Q8.0 input
    output reg [9:0] out // Q6.4 output
);

    always @(*) begin
        casez (in)
            8'd0  : out = 10'd0;   // 0^0.70 ~= 0.000000
            8'd1  : out = 10'd16;  // 1^0.70 ~= 1.000000
            8'd2  : out = 10'd26;  // 2^0.70 ~= 1.624505
            8'd3  : out = 10'd35;  // 3^0.70 ~= 2.157669
            8'd4  : out = 10'd42;  // 4^0.70 ~= 2.639016
            8'd5  : out = 10'd49;  // 5^0.70 ~= 3.085169
            8'd6  : out = 10'd56;  // 6^0.70 ~= 3.505144
            8'd7  : out = 10'd62;  // 7^0.70 ~= 3.904529
            8'd8  : out = 10'd69;  // 8^0.70 ~= 4.287094
            8'd9  : out = 10'd74;  // 9^0.70 ~= 4.655537
            8'd10 : out = 10'd80;  // 10^0.70 ~= 5.011872
            8'd11 : out = 10'd86;  // 11^0.70 ~= 5.357657
            8'd12 : out = 10'd91;  // 12^0.70 ~= 5.694123
            8'd13 : out = 10'd96;  // 13^0.70 ~= 6.022272
            8'd14 : out = 10'd101;  // 14^0.70 ~= 6.342926
            8'd15 : out = 10'd107;  // 15^0.70 ~= 6.656775
            8'd16 : out = 10'd111;  // 16^0.70 ~= 6.964405
            8'd17 : out = 10'd116;  // 17^0.70 ~= 7.266315
            8'd18 : out = 10'd121;  // 18^0.70 ~= 7.562942
            8'd19 : out = 10'd126;  // 19^0.70 ~= 7.854662
            8'd20 : out = 10'd130;  // 20^0.70 ~= 8.141811
            8'd21 : out = 10'd135;  // 21^0.70 ~= 8.424682
            8'd22 : out = 10'd139;  // 22^0.70 ~= 8.703539
            8'd23 : out = 10'd144;  // 23^0.70 ~= 8.978618
            8'd24 : out = 10'd148;  // 24^0.70 ~= 9.250131
            8'd25 : out = 10'd152;  // 25^0.70 ~= 9.518270
            8'd26 : out = 10'd157;  // 26^0.70 ~= 9.783209
            8'd27 : out = 10'd161;  // 27^0.70 ~= 10.045109
            8'd28 : out = 10'd165;  // 28^0.70 ~= 10.304113
            8'd29 : out = 10'd169;  // 29^0.70 ~= 10.560357
            8'd30 : out = 10'd173;  // 30^0.70 ~= 10.813963
            8'd31 : out = 10'd177;  // 31^0.70 ~= 11.065045
            8'd32 : out = 10'd181;  // 32^0.70 ~= 11.313708
            8'd33 : out = 10'd185;  // 33^0.70 ~= 11.560051
            8'd34 : out = 10'd189;  // 34^0.70 ~= 11.804164
            8'd35 : out = 10'd193;  // 35^0.70 ~= 12.046132
            8'd36 : out = 10'd197;  // 36^0.70 ~= 12.286035
            8'd37 : out = 10'd200;  // 37^0.70 ~= 12.523947
            8'd38 : out = 10'd204;  // 38^0.70 ~= 12.759937
            8'd39 : out = 10'd208;  // 39^0.70 ~= 12.994071
            8'd40 : out = 10'd212;  // 40^0.70 ~= 13.226410
            8'd41 : out = 10'd215;  // 41^0.70 ~= 13.457014
            8'd42 : out = 10'd219;  // 42^0.70 ~= 13.685936
            8'd43 : out = 10'd223;  // 43^0.70 ~= 13.913229
            8'd44 : out = 10'd226;  // 44^0.70 ~= 14.138941
            8'd45 : out = 10'd230;  // 45^0.70 ~= 14.363119
            8'd46 : out = 10'd233;  // 46^0.70 ~= 14.585808
            8'd47 : out = 10'd237;  // 47^0.70 ~= 14.807049
            8'd48 : out = 10'd240;  // 48^0.70 ~= 15.026882
            8'd49 : out = 10'd244;  // 49^0.70 ~= 15.245345
            8'd50 : out = 10'd247;  // 50^0.70 ~= 15.462475
            8'd51 : out = 10'd251;  // 51^0.70 ~= 15.678306
            8'd52 : out = 10'd254;  // 52^0.70 ~= 15.892870
            8'd53 : out = 10'd258;  // 53^0.70 ~= 16.106201
            8'd54 : out = 10'd261;  // 54^0.70 ~= 16.318327
            8'd55 : out = 10'd264;  // 55^0.70 ~= 16.529278
            8'd56 : out = 10'd268;  // 56^0.70 ~= 16.739081
            8'd57 : out = 10'd271;  // 57^0.70 ~= 16.947764
            8'd58 : out = 10'd274;  // 58^0.70 ~= 17.155350
            8'd59 : out = 10'd278;  // 59^0.70 ~= 17.361866
            8'd60 : out = 10'd281;  // 60^0.70 ~= 17.567335
            8'd61 : out = 10'd284;  // 61^0.70 ~= 17.771778
            8'd62 : out = 10'd288;  // 62^0.70 ~= 17.975219
            8'd63 : out = 10'd291;  // 63^0.70 ~= 18.177677
            8'd64 : out = 10'd294;  // 64^0.70 ~= 18.379174
            8'd65 : out = 10'd297;  // 65^0.70 ~= 18.579728
            8'd66 : out = 10'd300;  // 66^0.70 ~= 18.779359
            8'd67 : out = 10'd304;  // 67^0.70 ~= 18.978084
            8'd68 : out = 10'd307;  // 68^0.70 ~= 19.175921
            8'd69 : out = 10'd310;  // 69^0.70 ~= 19.372888
            8'd70 : out = 10'd313;  // 70^0.70 ~= 19.569000
            8'd71 : out = 10'd316;  // 71^0.70 ~= 19.764273
            8'd72 : out = 10'd319;  // 72^0.70 ~= 19.958723
            8'd73 : out = 10'd322;  // 73^0.70 ~= 20.152364
            8'd74 : out = 10'd326;  // 74^0.70 ~= 20.345211
            8'd75 : out = 10'd329;  // 75^0.70 ~= 20.537278
            8'd76 : out = 10'd332;  // 76^0.70 ~= 20.728578
            8'd77 : out = 10'd335;  // 77^0.70 ~= 20.919125
            8'd78 : out = 10'd338;  // 78^0.70 ~= 21.108930
            8'd79 : out = 10'd341;  // 79^0.70 ~= 21.298007
            8'd80 : out = 10'd344;  // 80^0.70 ~= 21.486367
            8'd81 : out = 10'd347;  // 81^0.70 ~= 21.674022
            8'd82 : out = 10'd350;  // 82^0.70 ~= 21.860984
            8'd83 : out = 10'd353;  // 83^0.70 ~= 22.047262
            8'd84 : out = 10'd356;  // 84^0.70 ~= 22.232869
            8'd85 : out = 10'd359;  // 85^0.70 ~= 22.417813
            8'd86 : out = 10'd362;  // 86^0.70 ~= 22.602106
            8'd87 : out = 10'd365;  // 87^0.70 ~= 22.785758
            8'd88 : out = 10'd368;  // 88^0.70 ~= 22.968777
            8'd89 : out = 10'd370;  // 89^0.70 ~= 23.151173
            8'd90 : out = 10'd373;  // 90^0.70 ~= 23.332956
            8'd91 : out = 10'd376;  // 91^0.70 ~= 23.514133
            8'd92 : out = 10'd379;  // 92^0.70 ~= 23.694714
            8'd93 : out = 10'd382;  // 93^0.70 ~= 23.874708
            8'd94 : out = 10'd385;  // 94^0.70 ~= 24.054121
            8'd95 : out = 10'd388;  // 95^0.70 ~= 24.232963
            8'd96 : out = 10'd391;  // 96^0.70 ~= 24.411241
            8'd97 : out = 10'd393;  // 97^0.70 ~= 24.588963
            8'd98 : out = 10'd396;  // 98^0.70 ~= 24.766136
            8'd99 : out = 10'd399;  // 99^0.70 ~= 24.942767
            8'd100: out = 10'd402;  // 100^0.70 ~= 25.118864
            8'd101: out = 10'd405;  // 101^0.70 ~= 25.294434
            8'd102: out = 10'd408;  // 102^0.70 ~= 25.469482
            8'd103: out = 10'd410;  // 103^0.70 ~= 25.644017
            8'd104: out = 10'd413;  // 104^0.70 ~= 25.818044
            8'd105: out = 10'd416;  // 105^0.70 ~= 25.991570
            8'd106: out = 10'd419;  // 106^0.70 ~= 26.164600
            8'd107: out = 10'd421;  // 107^0.70 ~= 26.337142
            8'd108: out = 10'd424;  // 108^0.70 ~= 26.509200
            8'd109: out = 10'd427;  // 109^0.70 ~= 26.680782
            8'd110: out = 10'd430;  // 110^0.70 ~= 26.851891
            8'd111: out = 10'd432;  // 111^0.70 ~= 27.022535
            8'd112: out = 10'd435;  // 112^0.70 ~= 27.192718
            8'd113: out = 10'd438;  // 113^0.70 ~= 27.362446
            8'd114: out = 10'd441;  // 114^0.70 ~= 27.531723
            8'd115: out = 10'd443;  // 115^0.70 ~= 27.700556
            8'd116: out = 10'd446;  // 116^0.70 ~= 27.868949
            8'd117: out = 10'd449;  // 117^0.70 ~= 28.036907
            8'd118: out = 10'd451;  // 118^0.70 ~= 28.204435
            8'd119: out = 10'd454;  // 119^0.70 ~= 28.371538
            8'd120: out = 10'd457;  // 120^0.70 ~= 28.538219
            8'd121: out = 10'd459;  // 121^0.70 ~= 28.704485
            8'd122: out = 10'd462;  // 122^0.70 ~= 28.870339
            8'd123: out = 10'd465;  // 123^0.70 ~= 29.035785
            8'd124: out = 10'd467;  // 124^0.70 ~= 29.200829
            8'd125: out = 10'd470;  // 125^0.70 ~= 29.365474
            8'd126: out = 10'd472;  // 126^0.70 ~= 29.529724
            8'd127: out = 10'd475;  // 127^0.70 ~= 29.693583
            8'd128: out = 10'd478;  // 128^0.70 ~= 29.857056
            8'd129: out = 10'd480;  // 129^0.70 ~= 30.020146
            8'd130: out = 10'd483;  // 130^0.70 ~= 30.182857
            8'd131: out = 10'd486;  // 131^0.70 ~= 30.345193
            8'd132: out = 10'd488;  // 132^0.70 ~= 30.507158
            8'd133: out = 10'd491;  // 133^0.70 ~= 30.668755
            8'd134: out = 10'd493;  // 134^0.70 ~= 30.829988
            8'd135: out = 10'd496;  // 135^0.70 ~= 30.990861
            8'd136: out = 10'd498;  // 136^0.70 ~= 31.151376
            8'd137: out = 10'd501;  // 137^0.70 ~= 31.311538
            8'd138: out = 10'd504;  // 138^0.70 ~= 31.471349
            8'd139: out = 10'd506;  // 139^0.70 ~= 31.630813
            8'd140: out = 10'd509;  // 140^0.70 ~= 31.789934
            8'd141: out = 10'd511;  // 141^0.70 ~= 31.948714
            8'd142: out = 10'd514;  // 142^0.70 ~= 32.107156
            8'd143: out = 10'd516;  // 143^0.70 ~= 32.265264
            8'd144: out = 10'd519;  // 144^0.70 ~= 32.423041
            8'd145: out = 10'd521;  // 145^0.70 ~= 32.580489
            8'd146: out = 10'd524;  // 146^0.70 ~= 32.737612
            8'd147: out = 10'd526;  // 147^0.70 ~= 32.894413
            8'd148: out = 10'd529;  // 148^0.70 ~= 33.050893
            8'd149: out = 10'd531;  // 149^0.70 ~= 33.207057
            8'd150: out = 10'd534;  // 150^0.70 ~= 33.362907
            8'd151: out = 10'd536;  // 151^0.70 ~= 33.518445
            8'd152: out = 10'd539;  // 152^0.70 ~= 33.673675
            8'd153: out = 10'd541;  // 153^0.70 ~= 33.828598
            8'd154: out = 10'd544;  // 154^0.70 ~= 33.983218
            8'd155: out = 10'd546;  // 155^0.70 ~= 34.137537
            8'd156: out = 10'd549;  // 156^0.70 ~= 34.291558
            8'd157: out = 10'd551;  // 157^0.70 ~= 34.445283
            8'd158: out = 10'd554;  // 158^0.70 ~= 34.598714
            8'd159: out = 10'd556;  // 159^0.70 ~= 34.751855
            8'd160: out = 10'd558;  // 160^0.70 ~= 34.904706
            8'd161: out = 10'd561;  // 161^0.70 ~= 35.057272
            8'd162: out = 10'd563;  // 162^0.70 ~= 35.209553
            8'd163: out = 10'd566;  // 163^0.70 ~= 35.361552
            8'd164: out = 10'd568;  // 164^0.70 ~= 35.513272
            8'd165: out = 10'd571;  // 165^0.70 ~= 35.664715
            8'd166: out = 10'd573;  // 166^0.70 ~= 35.815883
            8'd167: out = 10'd575;  // 167^0.70 ~= 35.966778
            8'd168: out = 10'd578;  // 168^0.70 ~= 36.117402
            8'd169: out = 10'd580;  // 169^0.70 ~= 36.267757
            8'd170: out = 10'd583;  // 170^0.70 ~= 36.417845
            8'd171: out = 10'd585;  // 171^0.70 ~= 36.567669
            8'd172: out = 10'd587;  // 172^0.70 ~= 36.717230
            8'd173: out = 10'd590;  // 173^0.70 ~= 36.866531
            8'd174: out = 10'd592;  // 174^0.70 ~= 37.015573
            8'd175: out = 10'd595;  // 175^0.70 ~= 37.164358
            8'd176: out = 10'd597;  // 176^0.70 ~= 37.312888
            8'd177: out = 10'd599;  // 177^0.70 ~= 37.461166
            8'd178: out = 10'd602;  // 178^0.70 ~= 37.609192
            8'd179: out = 10'd604;  // 179^0.70 ~= 37.756969
            8'd180: out = 10'd606;  // 180^0.70 ~= 37.904498
            8'd181: out = 10'd609;  // 181^0.70 ~= 38.051782
            8'd182: out = 10'd611;  // 182^0.70 ~= 38.198822
            8'd183: out = 10'd614;  // 183^0.70 ~= 38.345620
            8'd184: out = 10'd616;  // 184^0.70 ~= 38.492177
            8'd185: out = 10'd618;  // 185^0.70 ~= 38.638496
            8'd186: out = 10'd621;  // 186^0.70 ~= 38.784577
            8'd187: out = 10'd623;  // 187^0.70 ~= 38.930423
            8'd188: out = 10'd625;  // 188^0.70 ~= 39.076035
            8'd189: out = 10'd628;  // 189^0.70 ~= 39.221415
            8'd190: out = 10'd630;  // 190^0.70 ~= 39.366565
            8'd191: out = 10'd632;  // 191^0.70 ~= 39.511485
            8'd192: out = 10'd634;  // 192^0.70 ~= 39.656178
            8'd193: out = 10'd637;  // 193^0.70 ~= 39.800646
            8'd194: out = 10'd639;  // 194^0.70 ~= 39.944888
            8'd195: out = 10'd641;  // 195^0.70 ~= 40.088908
            8'd196: out = 10'd644;  // 196^0.70 ~= 40.232707
            8'd197: out = 10'd646;  // 197^0.70 ~= 40.376285
            8'd198: out = 10'd648;  // 198^0.70 ~= 40.519645
            8'd199: out = 10'd651;  // 199^0.70 ~= 40.662788
            8'd200: out = 10'd653;  // 200^0.70 ~= 40.805715
            8'd201: out = 10'd655;  // 201^0.70 ~= 40.948429
            8'd202: out = 10'd657;  // 202^0.70 ~= 41.090929
            8'd203: out = 10'd660;  // 203^0.70 ~= 41.233218
            8'd204: out = 10'd662;  // 204^0.70 ~= 41.375296
            8'd205: out = 10'd664;  // 205^0.70 ~= 41.517166
            8'd206: out = 10'd667;  // 206^0.70 ~= 41.658829
            8'd207: out = 10'd669;  // 207^0.70 ~= 41.800285
            8'd208: out = 10'd671;  // 208^0.70 ~= 41.941536
            8'd209: out = 10'd673;  // 209^0.70 ~= 42.082584
            8'd210: out = 10'd676;  // 210^0.70 ~= 42.223430
            8'd211: out = 10'd678;  // 211^0.70 ~= 42.364074
            8'd212: out = 10'd680;  // 212^0.70 ~= 42.504519
            8'd213: out = 10'd682;  // 213^0.70 ~= 42.644765
            8'd214: out = 10'd685;  // 214^0.70 ~= 42.784813
            8'd215: out = 10'd687;  // 215^0.70 ~= 42.924666
            8'd216: out = 10'd689;  // 216^0.70 ~= 43.064323
            8'd217: out = 10'd691;  // 217^0.70 ~= 43.203787
            8'd218: out = 10'd693;  // 218^0.70 ~= 43.343058
            8'd219: out = 10'd696;  // 219^0.70 ~= 43.482137
            8'd220: out = 10'd698;  // 220^0.70 ~= 43.621026
            8'd221: out = 10'd700;  // 221^0.70 ~= 43.759726
            8'd222: out = 10'd702;  // 222^0.70 ~= 43.898237
            8'd223: out = 10'd705;  // 223^0.70 ~= 44.036562
            8'd224: out = 10'd707;  // 224^0.70 ~= 44.174700
            8'd225: out = 10'd709;  // 225^0.70 ~= 44.312654
            8'd226: out = 10'd711;  // 226^0.70 ~= 44.450424
            8'd227: out = 10'd713;  // 227^0.70 ~= 44.588011
            8'd228: out = 10'd716;  // 228^0.70 ~= 44.725416
            8'd229: out = 10'd718;  // 229^0.70 ~= 44.862641
            8'd230: out = 10'd720;  // 230^0.70 ~= 44.999686
            8'd231: out = 10'd722;  // 231^0.70 ~= 45.136553
            8'd232: out = 10'd724;  // 232^0.70 ~= 45.273241
            8'd233: out = 10'd727;  // 233^0.70 ~= 45.409754
            8'd234: out = 10'd729;  // 234^0.70 ~= 45.546090
            8'd235: out = 10'd731;  // 235^0.70 ~= 45.682252
            8'd236: out = 10'd733;  // 236^0.70 ~= 45.818240
            8'd237: out = 10'd735;  // 237^0.70 ~= 45.954055
            8'd238: out = 10'd737;  // 238^0.70 ~= 46.089699
            8'd239: out = 10'd740;  // 239^0.70 ~= 46.225171
            8'd240: out = 10'd742;  // 240^0.70 ~= 46.360474
            8'd241: out = 10'd744;  // 241^0.70 ~= 46.495608
            8'd242: out = 10'd746;  // 242^0.70 ~= 46.630573
            8'd243: out = 10'd748;  // 243^0.70 ~= 46.765372
            8'd244: out = 10'd750;  // 244^0.70 ~= 46.900004
            8'd245: out = 10'd753;  // 245^0.70 ~= 47.034470
            8'd246: out = 10'd755;  // 246^0.70 ~= 47.168773
            8'd247: out = 10'd757;  // 247^0.70 ~= 47.302911
            8'd248: out = 10'd759;  // 248^0.70 ~= 47.436887
            8'd249: out = 10'd761;  // 249^0.70 ~= 47.570700
            8'd250: out = 10'd763;  // 250^0.70 ~= 47.704353
            8'd251: out = 10'd765;  // 251^0.70 ~= 47.837845
            8'd252: out = 10'd768;  // 252^0.70 ~= 47.971177
            8'd253: out = 10'd770;  // 253^0.70 ~= 48.104352
            8'd254: out = 10'd772;  // 254^0.70 ~= 48.237368
            8'd255: out = 10'd774;  // 255^0.70 ~= 48.370227
            default: out = 10'd0;
        endcase
    end
endmodule
