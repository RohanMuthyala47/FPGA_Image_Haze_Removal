// Compute ω * Pc / Ac
module Multiplier_TE (
    input         clk,
    input         rst,
    
    input  [7:0]  Fc,     // Filter result
    input  [13:0] Inv_Ac, // Scaled Inverted Atmospheric Light value in Q0.12 format (ω * 1/Ac) 
    
    output [7:0] product // ω * min(Pc / Ac) ; c ∈ {R, G, B} in Q0.8 format
);
    
    // Pipeline registers
    reg [17:0] result_P;
    
    // Pipeline inputs to reduce fan-out
    always @(posedge clk) begin
        if(rst) begin
            result_P <= 0;
        end
        else begin
            result_P <= Fc * Inv_Ac[13:4]; // Q8.10
        end
    end
    
    assign product = result_P[9:2]; // Scale down to Q0.8 and eliminate overflow
    
endmodule
