module Trans_LUT (
    input      [15:0] x, // Q0.16 Transmission value input (unsigned)
    output reg [15:0] y  // Q2.14 Inverse Transmission value output (unsigned)
);
    
    always @(*) begin
        casez(x[15:4])
            12'd   0: y = 16'h4000;
            12'd   1: y = 16'hFFFF;
            12'd   2: y = 16'hFFFF;
            12'd   3: y = 16'hFFFF;
            12'd   4: y = 16'hFFFF;
            12'd   5: y = 16'hFFFF;
            12'd   6: y = 16'hFFFF;
            12'd   7: y = 16'hFFFF;
            12'd   8: y = 16'hFFFF;
            12'd   9: y = 16'hFFFF;
            12'd  10: y = 16'hFFFF;
            12'd  11: y = 16'hFFFF;
            12'd  12: y = 16'hFFFF;
            12'd  13: y = 16'hFFFF;
            12'd  14: y = 16'hFFFF;
            12'd  15: y = 16'hFFFF;
            12'd  16: y = 16'hFFFF;
            12'd  17: y = 16'hFFFF;
            12'd  18: y = 16'hFFFF;
            12'd  19: y = 16'hFFFF;
            12'd  20: y = 16'hFFFF;
            12'd  21: y = 16'hFFFF;
            12'd  22: y = 16'hFFFF;
            12'd  23: y = 16'hFFFF;
            12'd  24: y = 16'hFFFF;
            12'd  25: y = 16'hFFFF;
            12'd  26: y = 16'hFFFF;
            12'd  27: y = 16'hFFFF;
            12'd  28: y = 16'hFFFF;
            12'd  29: y = 16'hFFFF;
            12'd  30: y = 16'hFFFF;
            12'd  31: y = 16'hFFFF;
            12'd  32: y = 16'hFFFF;
            12'd  33: y = 16'hFFFF;
            12'd  34: y = 16'hFFFF;
            12'd  35: y = 16'hFFFF;
            12'd  36: y = 16'hFFFF;
            12'd  37: y = 16'hFFFF;
            12'd  38: y = 16'hFFFF;
            12'd  39: y = 16'hFFFF;
            12'd  40: y = 16'hFFFF;
            12'd  41: y = 16'hFFFF;
            12'd  42: y = 16'hFFFF;
            12'd  43: y = 16'hFFFF;
            12'd  44: y = 16'hFFFF;
            12'd  45: y = 16'hFFFF;
            12'd  46: y = 16'hFFFF;
            12'd  47: y = 16'hFFFF;
            12'd  48: y = 16'hFFFF;
            12'd  49: y = 16'hFFFF;
            12'd  50: y = 16'hFFFF;
            12'd  51: y = 16'hFFFF;
            12'd  52: y = 16'hFFFF;
            12'd  53: y = 16'hFFFF;
            12'd  54: y = 16'hFFFF;
            12'd  55: y = 16'hFFFF;
            12'd  56: y = 16'hFFFF;
            12'd  57: y = 16'hFFFF;
            12'd  58: y = 16'hFFFF;
            12'd  59: y = 16'hFFFF;
            12'd  60: y = 16'hFFFF;
            12'd  61: y = 16'hFFFF;
            12'd  62: y = 16'hFFFF;
            12'd  63: y = 16'hFFFF;
            12'd  64: y = 16'hFFFF;
            12'd  65: y = 16'hFFFF;
            12'd  66: y = 16'hFFFF;
            12'd  67: y = 16'hFFFF;
            12'd  68: y = 16'hFFFF;
            12'd  69: y = 16'hFFFF;
            12'd  70: y = 16'hFFFF;
            12'd  71: y = 16'hFFFF;
            12'd  72: y = 16'hFFFF;
            12'd  73: y = 16'hFFFF;
            12'd  74: y = 16'hFFFF;
            12'd  75: y = 16'hFFFF;
            12'd  76: y = 16'hFFFF;
            12'd  77: y = 16'hFFFF;
            12'd  78: y = 16'hFFFF;
            12'd  79: y = 16'hFFFF;
            12'd  80: y = 16'hFFFF;
            12'd  81: y = 16'hFFFF;
            12'd  82: y = 16'hFFFF;
            12'd  83: y = 16'hFFFF;
            12'd  84: y = 16'hFFFF;
            12'd  85: y = 16'hFFFF;
            12'd  86: y = 16'hFFFF;
            12'd  87: y = 16'hFFFF;
            12'd  88: y = 16'hFFFF;
            12'd  89: y = 16'hFFFF;
            12'd  90: y = 16'hFFFF;
            12'd  91: y = 16'hFFFF;
            12'd  92: y = 16'hFFFF;
            12'd  93: y = 16'hFFFF;
            12'd  94: y = 16'hFFFF;
            12'd  95: y = 16'hFFFF;
            12'd  96: y = 16'hFFFF;
            12'd  97: y = 16'hFFFF;
            12'd  98: y = 16'hFFFF;
            12'd  99: y = 16'hFFFF;
            12'd 100: y = 16'hFFFF;
            12'd 101: y = 16'hFFFF;
            12'd 102: y = 16'hFFFF;
            12'd 103: y = 16'hFFFF;
            12'd 104: y = 16'hFFFF;
            12'd 105: y = 16'hFFFF;
            12'd 106: y = 16'hFFFF;
            12'd 107: y = 16'hFFFF;
            12'd 108: y = 16'hFFFF;
            12'd 109: y = 16'hFFFF;
            12'd 110: y = 16'hFFFF;
            12'd 111: y = 16'hFFFF;
            12'd 112: y = 16'hFFFF;
            12'd 113: y = 16'hFFFF;
            12'd 114: y = 16'hFFFF;
            12'd 115: y = 16'hFFFF;
            12'd 116: y = 16'hFFFF;
            12'd 117: y = 16'hFFFF;
            12'd 118: y = 16'hFFFF;
            12'd 119: y = 16'hFFFF;
            12'd 120: y = 16'hFFFF;
            12'd 121: y = 16'hFFFF;
            12'd 122: y = 16'hFFFF;
            12'd 123: y = 16'hFFFF;
            12'd 124: y = 16'hFFFF;
            12'd 125: y = 16'hFFFF;
            12'd 126: y = 16'hFFFF;
            12'd 127: y = 16'hFFFF;
            12'd 128: y = 16'hFFFF;
            12'd 129: y = 16'hFFFF;
            12'd 130: y = 16'hFFFF;
            12'd 131: y = 16'hFFFF;
            12'd 132: y = 16'hFFFF;
            12'd 133: y = 16'hFFFF;
            12'd 134: y = 16'hFFFF;
            12'd 135: y = 16'hFFFF;
            12'd 136: y = 16'hFFFF;
            12'd 137: y = 16'hFFFF;
            12'd 138: y = 16'hFFFF;
            12'd 139: y = 16'hFFFF;
            12'd 140: y = 16'hFFFF;
            12'd 141: y = 16'hFFFF;
            12'd 142: y = 16'hFFFF;
            12'd 143: y = 16'hFFFF;
            12'd 144: y = 16'hFFFF;
            12'd 145: y = 16'hFFFF;
            12'd 146: y = 16'hFFFF;
            12'd 147: y = 16'hFFFF;
            12'd 148: y = 16'hFFFF;
            12'd 149: y = 16'hFFFF;
            12'd 150: y = 16'hFFFF;
            12'd 151: y = 16'hFFFF;
            12'd 152: y = 16'hFFFF;
            12'd 153: y = 16'hFFFF;
            12'd 154: y = 16'hFFFF;
            12'd 155: y = 16'hFFFF;
            12'd 156: y = 16'hFFFF;
            12'd 157: y = 16'hFFFF;
            12'd 158: y = 16'hFFFF;
            12'd 159: y = 16'hFFFF;
            12'd 160: y = 16'hFFFF;
            12'd 161: y = 16'hFFFF;
            12'd 162: y = 16'hFFFF;
            12'd 163: y = 16'hFFFF;
            12'd 164: y = 16'hFFFF;
            12'd 165: y = 16'hFFFF;
            12'd 166: y = 16'hFFFF;
            12'd 167: y = 16'hFFFF;
            12'd 168: y = 16'hFFFF;
            12'd 169: y = 16'hFFFF;
            12'd 170: y = 16'hFFFF;
            12'd 171: y = 16'hFFFF;
            12'd 172: y = 16'hFFFF;
            12'd 173: y = 16'hFFFF;
            12'd 174: y = 16'hFFFF;
            12'd 175: y = 16'hFFFF;
            12'd 176: y = 16'hFFFF;
            12'd 177: y = 16'hFFFF;
            12'd 178: y = 16'hFFFF;
            12'd 179: y = 16'hFFFF;
            12'd 180: y = 16'hFFFF;
            12'd 181: y = 16'hFFFF;
            12'd 182: y = 16'hFFFF;
            12'd 183: y = 16'hFFFF;
            12'd 184: y = 16'hFFFF;
            12'd 185: y = 16'hFFFF;
            12'd 186: y = 16'hFFFF;
            12'd 187: y = 16'hFFFF;
            12'd 188: y = 16'hFFFF;
            12'd 189: y = 16'hFFFF;
            12'd 190: y = 16'hFFFF;
            12'd 191: y = 16'hFFFF;
            12'd 192: y = 16'hFFFF;
            12'd 193: y = 16'hFFFF;
            12'd 194: y = 16'hFFFF;
            12'd 195: y = 16'hFFFF;
            12'd 196: y = 16'hFFFF;
            12'd 197: y = 16'hFFFF;
            12'd 198: y = 16'hFFFF;
            12'd 199: y = 16'hFFFF;
            12'd 200: y = 16'hFFFF;
            12'd 201: y = 16'hFFFF;
            12'd 202: y = 16'hFFFF;
            12'd 203: y = 16'hFFFF;
            12'd 204: y = 16'hFFFF;
            12'd 205: y = 16'hFFFF;
            12'd 206: y = 16'hFFFF;
            12'd 207: y = 16'hFFFF;
            12'd 208: y = 16'hFFFF;
            12'd 209: y = 16'hFFFF;
            12'd 210: y = 16'hFFFF;
            12'd 211: y = 16'hFFFF;
            12'd 212: y = 16'hFFFF;
            12'd 213: y = 16'hFFFF;
            12'd 214: y = 16'hFFFF;
            12'd 215: y = 16'hFFFF;
            12'd 216: y = 16'hFFFF;
            12'd 217: y = 16'hFFFF;
            12'd 218: y = 16'hFFFF;
            12'd 219: y = 16'hFFFF;
            12'd 220: y = 16'hFFFF;
            12'd 221: y = 16'hFFFF;
            12'd 222: y = 16'hFFFF;
            12'd 223: y = 16'hFFFF;
            12'd 224: y = 16'hFFFF;
            12'd 225: y = 16'hFFFF;
            12'd 226: y = 16'hFFFF;
            12'd 227: y = 16'hFFFF;
            12'd 228: y = 16'hFFFF;
            12'd 229: y = 16'hFFFF;
            12'd 230: y = 16'hFFFF;
            12'd 231: y = 16'hFFFF;
            12'd 232: y = 16'hFFFF;
            12'd 233: y = 16'hFFFF;
            12'd 234: y = 16'hFFFF;
            12'd 235: y = 16'hFFFF;
            12'd 236: y = 16'hFFFF;
            12'd 237: y = 16'hFFFF;
            12'd 238: y = 16'hFFFF;
            12'd 239: y = 16'hFFFF;
            12'd 240: y = 16'hFFFF;
            12'd 241: y = 16'hFFFF;
            12'd 242: y = 16'hFFFF;
            12'd 243: y = 16'hFFFF;
            12'd 244: y = 16'hFFFF;
            12'd 245: y = 16'hFFFF;
            12'd 246: y = 16'hFFFF;
            12'd 247: y = 16'hFFFF;
            12'd 248: y = 16'hFFFF;
            12'd 249: y = 16'hFFFF;
            12'd 250: y = 16'hFFFF;
            12'd 251: y = 16'hFFFF;
            12'd 252: y = 16'hFFFF;
            12'd 253: y = 16'hFFFF;
            12'd 254: y = 16'hFFFF;
            12'd 255: y = 16'hFFFF;
            12'd 256: y = 16'hFFFF;
            12'd 257: y = 16'hFFFF;
            12'd 258: y = 16'hFFFF;
            12'd 259: y = 16'hFFFF;
            12'd 260: y = 16'hFFFF;
            12'd 261: y = 16'hFFFF;
            12'd 262: y = 16'hFFFF;
            12'd 263: y = 16'hFFFF;
            12'd 264: y = 16'hFFFF;
            12'd 265: y = 16'hFFFF;
            12'd 266: y = 16'hFFFF;
            12'd 267: y = 16'hFFFF;
            12'd 268: y = 16'hFFFF;
            12'd 269: y = 16'hFFFF;
            12'd 270: y = 16'hFFFF;
            12'd 271: y = 16'hFFFF;
            12'd 272: y = 16'hFFFF;
            12'd 273: y = 16'hFFFF;
            12'd 274: y = 16'hFFFF;
            12'd 275: y = 16'hFFFF;
            12'd 276: y = 16'hFFFF;
            12'd 277: y = 16'hFFFF;
            12'd 278: y = 16'hFFFF;
            12'd 279: y = 16'hFFFF;
            12'd 280: y = 16'hFFFF;
            12'd 281: y = 16'hFFFF;
            12'd 282: y = 16'hFFFF;
            12'd 283: y = 16'hFFFF;
            12'd 284: y = 16'hFFFF;
            12'd 285: y = 16'hFFFF;
            12'd 286: y = 16'hFFFF;
            12'd 287: y = 16'hFFFF;
            12'd 288: y = 16'hFFFF;
            12'd 289: y = 16'hFFFF;
            12'd 290: y = 16'hFFFF;
            12'd 291: y = 16'hFFFF;
            12'd 292: y = 16'hFFFF;
            12'd 293: y = 16'hFFFF;
            12'd 294: y = 16'hFFFF;
            12'd 295: y = 16'hFFFF;
            12'd 296: y = 16'hFFFF;
            12'd 297: y = 16'hFFFF;
            12'd 298: y = 16'hFFFF;
            12'd 299: y = 16'hFFFF;
            12'd 300: y = 16'hFFFF;
            12'd 301: y = 16'hFFFF;
            12'd 302: y = 16'hFFFF;
            12'd 303: y = 16'hFFFF;
            12'd 304: y = 16'hFFFF;
            12'd 305: y = 16'hFFFF;
            12'd 306: y = 16'hFFFF;
            12'd 307: y = 16'hFFFF;
            12'd 308: y = 16'hFFFF;
            12'd 309: y = 16'hFFFF;
            12'd 310: y = 16'hFFFF;
            12'd 311: y = 16'hFFFF;
            12'd 312: y = 16'hFFFF;
            12'd 313: y = 16'hFFFF;
            12'd 314: y = 16'hFFFF;
            12'd 315: y = 16'hFFFF;
            12'd 316: y = 16'hFFFF;
            12'd 317: y = 16'hFFFF;
            12'd 318: y = 16'hFFFF;
            12'd 319: y = 16'hFFFF;
            12'd 320: y = 16'hFFFF;
            12'd 321: y = 16'hFFFF;
            12'd 322: y = 16'hFFFF;
            12'd 323: y = 16'hFFFF;
            12'd 324: y = 16'hFFFF;
            12'd 325: y = 16'hFFFF;
            12'd 326: y = 16'hFFFF;
            12'd 327: y = 16'hFFFF;
            12'd 328: y = 16'hFFFF;
            12'd 329: y = 16'hFFFF;
            12'd 330: y = 16'hFFFF;
            12'd 331: y = 16'hFFFF;
            12'd 332: y = 16'hFFFF;
            12'd 333: y = 16'hFFFF;
            12'd 334: y = 16'hFFFF;
            12'd 335: y = 16'hFFFF;
            12'd 336: y = 16'hFFFF;
            12'd 337: y = 16'hFFFF;
            12'd 338: y = 16'hFFFF;
            12'd 339: y = 16'hFFFF;
            12'd 340: y = 16'hFFFF;
            12'd 341: y = 16'hFFFF;
            12'd 342: y = 16'hFFFF;
            12'd 343: y = 16'hFFFF;
            12'd 344: y = 16'hFFFF;
            12'd 345: y = 16'hFFFF;
            12'd 346: y = 16'hFFFF;
            12'd 347: y = 16'hFFFF;
            12'd 348: y = 16'hFFFF;
            12'd 349: y = 16'hFFFF;
            12'd 350: y = 16'hFFFF;
            12'd 351: y = 16'hFFFF;
            12'd 352: y = 16'hFFFF;
            12'd 353: y = 16'hFFFF;
            12'd 354: y = 16'hFFFF;
            12'd 355: y = 16'hFFFF;
            12'd 356: y = 16'hFFFF;
            12'd 357: y = 16'hFFFF;
            12'd 358: y = 16'hFFFF;
            12'd 359: y = 16'hFFFF;
            12'd 360: y = 16'hFFFF;
            12'd 361: y = 16'hFFFF;
            12'd 362: y = 16'hFFFF;
            12'd 363: y = 16'hFFFF;
            12'd 364: y = 16'hFFFF;
            12'd 365: y = 16'hFFFF;
            12'd 366: y = 16'hFFFF;
            12'd 367: y = 16'hFFFF;
            12'd 368: y = 16'hFFFF;
            12'd 369: y = 16'hFFFF;
            12'd 370: y = 16'hFFFF;
            12'd 371: y = 16'hFFFF;
            12'd 372: y = 16'hFFFF;
            12'd 373: y = 16'hFFFF;
            12'd 374: y = 16'hFFFF;
            12'd 375: y = 16'hFFFF;
            12'd 376: y = 16'hFFFF;
            12'd 377: y = 16'hFFFF;
            12'd 378: y = 16'hFFFF;
            12'd 379: y = 16'hFFFF;
            12'd 380: y = 16'hFFFF;
            12'd 381: y = 16'hFFFF;
            12'd 382: y = 16'hFFFF;
            12'd 383: y = 16'hFFFF;
            12'd 384: y = 16'hFFFF;
            12'd 385: y = 16'hFFFF;
            12'd 386: y = 16'hFFFF;
            12'd 387: y = 16'hFFFF;
            12'd 388: y = 16'hFFFF;
            12'd 389: y = 16'hFFFF;
            12'd 390: y = 16'hFFFF;
            12'd 391: y = 16'hFFFF;
            12'd 392: y = 16'hFFFF;
            12'd 393: y = 16'hFFFF;
            12'd 394: y = 16'hFFFF;
            12'd 395: y = 16'hFFFF;
            12'd 396: y = 16'hFFFF;
            12'd 397: y = 16'hFFFF;
            12'd 398: y = 16'hFFFF;
            12'd 399: y = 16'hFFFF;
            12'd 400: y = 16'hFFFF;
            12'd 401: y = 16'hFFFF;
            12'd 402: y = 16'hFFFF;
            12'd 403: y = 16'hFFFF;
            12'd 404: y = 16'hFFFF;
            12'd 405: y = 16'hFFFF;
            12'd 406: y = 16'hFFFF;
            12'd 407: y = 16'hFFFF;
            12'd 408: y = 16'hFFFF;
            12'd 409: y = 16'hFFFF;
            12'd 410: y = 16'hFFFF;
            12'd 411: y = 16'hFFFF;
            12'd 412: y = 16'hFFFF;
            12'd 413: y = 16'hFFFF;
            12'd 414: y = 16'hFFFF;
            12'd 415: y = 16'hFFFF;
            12'd 416: y = 16'hFFFF;
            12'd 417: y = 16'hFFFF;
            12'd 418: y = 16'hFFFF;
            12'd 419: y = 16'hFFFF;
            12'd 420: y = 16'hFFFF;
            12'd 421: y = 16'hFFFF;
            12'd 422: y = 16'hFFFF;
            12'd 423: y = 16'hFFFF;
            12'd 424: y = 16'hFFFF;
            12'd 425: y = 16'hFFFF;
            12'd 426: y = 16'hFFFF;
            12'd 427: y = 16'hFFFF;
            12'd 428: y = 16'hFFFF;
            12'd 429: y = 16'hFFFF;
            12'd 430: y = 16'hFFFF;
            12'd 431: y = 16'hFFFF;
            12'd 432: y = 16'hFFFF;
            12'd 433: y = 16'hFFFF;
            12'd 434: y = 16'hFFFF;
            12'd 435: y = 16'hFFFF;
            12'd 436: y = 16'hFFFF;
            12'd 437: y = 16'hFFFF;
            12'd 438: y = 16'hFFFF;
            12'd 439: y = 16'hFFFF;
            12'd 440: y = 16'hFFFF;
            12'd 441: y = 16'hFFFF;
            12'd 442: y = 16'hFFFF;
            12'd 443: y = 16'hFFFF;
            12'd 444: y = 16'hFFFF;
            12'd 445: y = 16'hFFFF;
            12'd 446: y = 16'hFFFF;
            12'd 447: y = 16'hFFFF;
            12'd 448: y = 16'hFFFF;
            12'd 449: y = 16'hFFFF;
            12'd 450: y = 16'hFFFF;
            12'd 451: y = 16'hFFFF;
            12'd 452: y = 16'hFFFF;
            12'd 453: y = 16'hFFFF;
            12'd 454: y = 16'hFFFF;
            12'd 455: y = 16'hFFFF;
            12'd 456: y = 16'hFFFF;
            12'd 457: y = 16'hFFFF;
            12'd 458: y = 16'hFFFF;
            12'd 459: y = 16'hFFFF;
            12'd 460: y = 16'hFFFF;
            12'd 461: y = 16'hFFFF;
            12'd 462: y = 16'hFFFF;
            12'd 463: y = 16'hFFFF;
            12'd 464: y = 16'hFFFF;
            12'd 465: y = 16'hFFFF;
            12'd 466: y = 16'hFFFF;
            12'd 467: y = 16'hFFFF;
            12'd 468: y = 16'hFFFF;
            12'd 469: y = 16'hFFFF;
            12'd 470: y = 16'hFFFF;
            12'd 471: y = 16'hFFFF;
            12'd 472: y = 16'hFFFF;
            12'd 473: y = 16'hFFFF;
            12'd 474: y = 16'hFFFF;
            12'd 475: y = 16'hFFFF;
            12'd 476: y = 16'hFFFF;
            12'd 477: y = 16'hFFFF;
            12'd 478: y = 16'hFFFF;
            12'd 479: y = 16'hFFFF;
            12'd 480: y = 16'hFFFF;
            12'd 481: y = 16'hFFFF;
            12'd 482: y = 16'hFFFF;
            12'd 483: y = 16'hFFFF;
            12'd 484: y = 16'hFFFF;
            12'd 485: y = 16'hFFFF;
            12'd 486: y = 16'hFFFF;
            12'd 487: y = 16'hFFFF;
            12'd 488: y = 16'hFFFF;
            12'd 489: y = 16'hFFFF;
            12'd 490: y = 16'hFFFF;
            12'd 491: y = 16'hFFFF;
            12'd 492: y = 16'hFFFF;
            12'd 493: y = 16'hFFFF;
            12'd 494: y = 16'hFFFF;
            12'd 495: y = 16'hFFFF;
            12'd 496: y = 16'hFFFF;
            12'd 497: y = 16'hFFFF;
            12'd 498: y = 16'hFFFF;
            12'd 499: y = 16'hFFFF;
            12'd 500: y = 16'hFFFF;
            12'd 501: y = 16'hFFFF;
            12'd 502: y = 16'hFFFF;
            12'd 503: y = 16'hFFFF;
            12'd 504: y = 16'hFFFF;
            12'd 505: y = 16'hFFFF;
            12'd 506: y = 16'hFFFF;
            12'd 507: y = 16'hFFFF;
            12'd 508: y = 16'hFFFF;
            12'd 509: y = 16'hFFFF;
            12'd 510: y = 16'hFFFF;
            12'd 511: y = 16'hFFFF;
            12'd 512: y = 16'hFFFF;
            12'd 513: y = 16'hFFFF;
            12'd 514: y = 16'hFFFF;
            12'd 515: y = 16'hFFFF;
            12'd 516: y = 16'hFFFF;
            12'd 517: y = 16'hFFFF;
            12'd 518: y = 16'hFFFF;
            12'd 519: y = 16'hFFFF;
            12'd 520: y = 16'hFFFF;
            12'd 521: y = 16'hFFFF;
            12'd 522: y = 16'hFFFF;
            12'd 523: y = 16'hFFFF;
            12'd 524: y = 16'hFFFF;
            12'd 525: y = 16'hFFFF;
            12'd 526: y = 16'hFFFF;
            12'd 527: y = 16'hFFFF;
            12'd 528: y = 16'hFFFF;
            12'd 529: y = 16'hFFFF;
            12'd 530: y = 16'hFFFF;
            12'd 531: y = 16'hFFFF;
            12'd 532: y = 16'hFFFF;
            12'd 533: y = 16'hFFFF;
            12'd 534: y = 16'hFFFF;
            12'd 535: y = 16'hFFFF;
            12'd 536: y = 16'hFFFF;
            12'd 537: y = 16'hFFFF;
            12'd 538: y = 16'hFFFF;
            12'd 539: y = 16'hFFFF;
            12'd 540: y = 16'hFFFF;
            12'd 541: y = 16'hFFFF;
            12'd 542: y = 16'hFFFF;
            12'd 543: y = 16'hFFFF;
            12'd 544: y = 16'hFFFF;
            12'd 545: y = 16'hFFFF;
            12'd 546: y = 16'hFFFF;
            12'd 547: y = 16'hFFFF;
            12'd 548: y = 16'hFFFF;
            12'd 549: y = 16'hFFFF;
            12'd 550: y = 16'hFFFF;
            12'd 551: y = 16'hFFFF;
            12'd 552: y = 16'hFFFF;
            12'd 553: y = 16'hFFFF;
            12'd 554: y = 16'hFFFF;
            12'd 555: y = 16'hFFFF;
            12'd 556: y = 16'hFFFF;
            12'd 557: y = 16'hFFFF;
            12'd 558: y = 16'hFFFF;
            12'd 559: y = 16'hFFFF;
            12'd 560: y = 16'hFFFF;
            12'd 561: y = 16'hFFFF;
            12'd 562: y = 16'hFFFF;
            12'd 563: y = 16'hFFFF;
            12'd 564: y = 16'hFFFF;
            12'd 565: y = 16'hFFFF;
            12'd 566: y = 16'hFFFF;
            12'd 567: y = 16'hFFFF;
            12'd 568: y = 16'hFFFF;
            12'd 569: y = 16'hFFFF;
            12'd 570: y = 16'hFFFF;
            12'd 571: y = 16'hFFFF;
            12'd 572: y = 16'hFFFF;
            12'd 573: y = 16'hFFFF;
            12'd 574: y = 16'hFFFF;
            12'd 575: y = 16'hFFFF;
            12'd 576: y = 16'hFFFF;
            12'd 577: y = 16'hFFFF;
            12'd 578: y = 16'hFFFF;
            12'd 579: y = 16'hFFFF;
            12'd 580: y = 16'hFFFF;
            12'd 581: y = 16'hFFFF;
            12'd 582: y = 16'hFFFF;
            12'd 583: y = 16'hFFFF;
            12'd 584: y = 16'hFFFF;
            12'd 585: y = 16'hFFFF;
            12'd 586: y = 16'hFFFF;
            12'd 587: y = 16'hFFFF;
            12'd 588: y = 16'hFFFF;
            12'd 589: y = 16'hFFFF;
            12'd 590: y = 16'hFFFF;
            12'd 591: y = 16'hFFFF;
            12'd 592: y = 16'hFFFF;
            12'd 593: y = 16'hFFFF;
            12'd 594: y = 16'hFFFF;
            12'd 595: y = 16'hFFFF;
            12'd 596: y = 16'hFFFF;
            12'd 597: y = 16'hFFFF;
            12'd 598: y = 16'hFFFF;
            12'd 599: y = 16'hFFFF;
            12'd 600: y = 16'hFFFF;
            12'd 601: y = 16'hFFFF;
            12'd 602: y = 16'hFFFF;
            12'd 603: y = 16'hFFFF;
            12'd 604: y = 16'hFFFF;
            12'd 605: y = 16'hFFFF;
            12'd 606: y = 16'hFFFF;
            12'd 607: y = 16'hFFFF;
            12'd 608: y = 16'hFFFF;
            12'd 609: y = 16'hFFFF;
            12'd 610: y = 16'hFFFF;
            12'd 611: y = 16'hFFFF;
            12'd 612: y = 16'hFFFF;
            12'd 613: y = 16'hFFFF;
            12'd 614: y = 16'hFFFF;
            12'd 615: y = 16'hFFFF;
            12'd 616: y = 16'hFFFF;
            12'd 617: y = 16'hFFFF;
            12'd 618: y = 16'hFFFF;
            12'd 619: y = 16'hFFFF;
            12'd 620: y = 16'hFFFF;
            12'd 621: y = 16'hFFFF;
            12'd 622: y = 16'hFFFF;
            12'd 623: y = 16'hFFFF;
            12'd 624: y = 16'hFFFF;
            12'd 625: y = 16'hFFFF;
            12'd 626: y = 16'hFFFF;
            12'd 627: y = 16'hFFFF;
            12'd 628: y = 16'hFFFF;
            12'd 629: y = 16'hFFFF;
            12'd 630: y = 16'hFFFF;
            12'd 631: y = 16'hFFFF;
            12'd 632: y = 16'hFFFF;
            12'd 633: y = 16'hFFFF;
            12'd 634: y = 16'hFFFF;
            12'd 635: y = 16'hFFFF;
            12'd 636: y = 16'hFFFF;
            12'd 637: y = 16'hFFFF;
            12'd 638: y = 16'hFFFF;
            12'd 639: y = 16'hFFFF;
            12'd 640: y = 16'hFFFF;
            12'd 641: y = 16'hFFFF;
            12'd 642: y = 16'hFFFF;
            12'd 643: y = 16'hFFFF;
            12'd 644: y = 16'hFFFF;
            12'd 645: y = 16'hFFFF;
            12'd 646: y = 16'hFFFF;
            12'd 647: y = 16'hFFFF;
            12'd 648: y = 16'hFFFF;
            12'd 649: y = 16'hFFFF;
            12'd 650: y = 16'hFFFF;
            12'd 651: y = 16'hFFFF;
            12'd 652: y = 16'hFFFF;
            12'd 653: y = 16'hFFFF;
            12'd 654: y = 16'hFFFF;
            12'd 655: y = 16'hFFFF;
            12'd 656: y = 16'hFFFF;
            12'd 657: y = 16'hFFFF;
            12'd 658: y = 16'hFFFF;
            12'd 659: y = 16'hFFFF;
            12'd 660: y = 16'hFFFF;
            12'd 661: y = 16'hFFFF;
            12'd 662: y = 16'hFFFF;
            12'd 663: y = 16'hFFFF;
            12'd 664: y = 16'hFFFF;
            12'd 665: y = 16'hFFFF;
            12'd 666: y = 16'hFFFF;
            12'd 667: y = 16'hFFFF;
            12'd 668: y = 16'hFFFF;
            12'd 669: y = 16'hFFFF;
            12'd 670: y = 16'hFFFF;
            12'd 671: y = 16'hFFFF;
            12'd 672: y = 16'hFFFF;
            12'd 673: y = 16'hFFFF;
            12'd 674: y = 16'hFFFF;
            12'd 675: y = 16'hFFFF;
            12'd 676: y = 16'hFFFF;
            12'd 677: y = 16'hFFFF;
            12'd 678: y = 16'hFFFF;
            12'd 679: y = 16'hFFFF;
            12'd 680: y = 16'hFFFF;
            12'd 681: y = 16'hFFFF;
            12'd 682: y = 16'hFFFF;
            12'd 683: y = 16'hFFFF;
            12'd 684: y = 16'hFFFF;
            12'd 685: y = 16'hFFFF;
            12'd 686: y = 16'hFFFF;
            12'd 687: y = 16'hFFFF;
            12'd 688: y = 16'hFFFF;
            12'd 689: y = 16'hFFFF;
            12'd 690: y = 16'hFFFF;
            12'd 691: y = 16'hFFFF;
            12'd 692: y = 16'hFFFF;
            12'd 693: y = 16'hFFFF;
            12'd 694: y = 16'hFFFF;
            12'd 695: y = 16'hFFFF;
            12'd 696: y = 16'hFFFF;
            12'd 697: y = 16'hFFFF;
            12'd 698: y = 16'hFFFF;
            12'd 699: y = 16'hFFFF;
            12'd 700: y = 16'hFFFF;
            12'd 701: y = 16'hFFFF;
            12'd 702: y = 16'hFFFF;
            12'd 703: y = 16'hFFFF;
            12'd 704: y = 16'hFFFF;
            12'd 705: y = 16'hFFFF;
            12'd 706: y = 16'hFFFF;
            12'd 707: y = 16'hFFFF;
            12'd 708: y = 16'hFFFF;
            12'd 709: y = 16'hFFFF;
            12'd 710: y = 16'hFFFF;
            12'd 711: y = 16'hFFFF;
            12'd 712: y = 16'hFFFF;
            12'd 713: y = 16'hFFFF;
            12'd 714: y = 16'hFFFF;
            12'd 715: y = 16'hFFFF;
            12'd 716: y = 16'hFFFF;
            12'd 717: y = 16'hFFFF;
            12'd 718: y = 16'hFFFF;
            12'd 719: y = 16'hFFFF;
            12'd 720: y = 16'hFFFF;
            12'd 721: y = 16'hFFFF;
            12'd 722: y = 16'hFFFF;
            12'd 723: y = 16'hFFFF;
            12'd 724: y = 16'hFFFF;
            12'd 725: y = 16'hFFFF;
            12'd 726: y = 16'hFFFF;
            12'd 727: y = 16'hFFFF;
            12'd 728: y = 16'hFFFF;
            12'd 729: y = 16'hFFFF;
            12'd 730: y = 16'hFFFF;
            12'd 731: y = 16'hFFFF;
            12'd 732: y = 16'hFFFF;
            12'd 733: y = 16'hFFFF;
            12'd 734: y = 16'hFFFF;
            12'd 735: y = 16'hFFFF;
            12'd 736: y = 16'hFFFF;
            12'd 737: y = 16'hFFFF;
            12'd 738: y = 16'hFFFF;
            12'd 739: y = 16'hFFFF;
            12'd 740: y = 16'hFFFF;
            12'd 741: y = 16'hFFFF;
            12'd 742: y = 16'hFFFF;
            12'd 743: y = 16'hFFFF;
            12'd 744: y = 16'hFFFF;
            12'd 745: y = 16'hFFFF;
            12'd 746: y = 16'hFFFF;
            12'd 747: y = 16'hFFFF;
            12'd 748: y = 16'hFFFF;
            12'd 749: y = 16'hFFFF;
            12'd 750: y = 16'hFFFF;
            12'd 751: y = 16'hFFFF;
            12'd 752: y = 16'hFFFF;
            12'd 753: y = 16'hFFFF;
            12'd 754: y = 16'hFFFF;
            12'd 755: y = 16'hFFFF;
            12'd 756: y = 16'hFFFF;
            12'd 757: y = 16'hFFFF;
            12'd 758: y = 16'hFFFF;
            12'd 759: y = 16'hFFFF;
            12'd 760: y = 16'hFFFF;
            12'd 761: y = 16'hFFFF;
            12'd 762: y = 16'hFFFF;
            12'd 763: y = 16'hFFFF;
            12'd 764: y = 16'hFFFF;
            12'd 765: y = 16'hFFFF;
            12'd 766: y = 16'hFFFF;
            12'd 767: y = 16'hFFFF;
            12'd 768: y = 16'hFFFF;
            12'd 769: y = 16'hFFFF;
            12'd 770: y = 16'hFFFF;
            12'd 771: y = 16'hFFFF;
            12'd 772: y = 16'hFFFF;
            12'd 773: y = 16'hFFFF;
            12'd 774: y = 16'hFFFF;
            12'd 775: y = 16'hFFFF;
            12'd 776: y = 16'hFFFF;
            12'd 777: y = 16'hFFFF;
            12'd 778: y = 16'hFFFF;
            12'd 779: y = 16'hFFFF;
            12'd 780: y = 16'hFFFF;
            12'd 781: y = 16'hFFFF;
            12'd 782: y = 16'hFFFF;
            12'd 783: y = 16'hFFFF;
            12'd 784: y = 16'hFFFF;
            12'd 785: y = 16'hFFFF;
            12'd 786: y = 16'hFFFF;
            12'd 787: y = 16'hFFFF;
            12'd 788: y = 16'hFFFF;
            12'd 789: y = 16'hFFFF;
            12'd 790: y = 16'hFFFF;
            12'd 791: y = 16'hFFFF;
            12'd 792: y = 16'hFFFF;
            12'd 793: y = 16'hFFFF;
            12'd 794: y = 16'hFFFF;
            12'd 795: y = 16'hFFFF;
            12'd 796: y = 16'hFFFF;
            12'd 797: y = 16'hFFFF;
            12'd 798: y = 16'hFFFF;
            12'd 799: y = 16'hFFFF;
            12'd 800: y = 16'hFFFF;
            12'd 801: y = 16'hFFFF;
            12'd 802: y = 16'hFFFF;
            12'd 803: y = 16'hFFFF;
            12'd 804: y = 16'hFFFF;
            12'd 805: y = 16'hFFFF;
            12'd 806: y = 16'hFFFF;
            12'd 807: y = 16'hFFFF;
            12'd 808: y = 16'hFFFF;
            12'd 809: y = 16'hFFFF;
            12'd 810: y = 16'hFFFF;
            12'd 811: y = 16'hFFFF;
            12'd 812: y = 16'hFFFF;
            12'd 813: y = 16'hFFFF;
            12'd 814: y = 16'hFFFF;
            12'd 815: y = 16'hFFFF;
            12'd 816: y = 16'hFFFF;
            12'd 817: y = 16'hFFFF;
            12'd 818: y = 16'hFFFF;
            12'd 819: y = 16'hFFFF;
            12'd 820: y = 16'hFFFF;
            12'd 821: y = 16'hFFFF;
            12'd 822: y = 16'hFFFF;
            12'd 823: y = 16'hFFFF;
            12'd 824: y = 16'hFFFF;
            12'd 825: y = 16'hFFFF;
            12'd 826: y = 16'hFFFF;
            12'd 827: y = 16'hFFFF;
            12'd 828: y = 16'hFFFF;
            12'd 829: y = 16'hFFFF;
            12'd 830: y = 16'hFFFF;
            12'd 831: y = 16'hFFFF;
            12'd 832: y = 16'hFFFF;
            12'd 833: y = 16'hFFFF;
            12'd 834: y = 16'hFFFF;
            12'd 835: y = 16'hFFFF;
            12'd 836: y = 16'hFFFF;
            12'd 837: y = 16'hFFFF;
            12'd 838: y = 16'hFFFF;
            12'd 839: y = 16'hFFFF;
            12'd 840: y = 16'hFFFF;
            12'd 841: y = 16'hFFFF;
            12'd 842: y = 16'hFFFF;
            12'd 843: y = 16'hFFFF;
            12'd 844: y = 16'hFFFF;
            12'd 845: y = 16'hFFFF;
            12'd 846: y = 16'hFFFF;
            12'd 847: y = 16'hFFFF;
            12'd 848: y = 16'hFFFF;
            12'd 849: y = 16'hFFFF;
            12'd 850: y = 16'hFFFF;
            12'd 851: y = 16'hFFFF;
            12'd 852: y = 16'hFFFF;
            12'd 853: y = 16'hFFFF;
            12'd 854: y = 16'hFFFF;
            12'd 855: y = 16'hFFFF;
            12'd 856: y = 16'hFFFF;
            12'd 857: y = 16'hFFFF;
            12'd 858: y = 16'hFFFF;
            12'd 859: y = 16'hFFFF;
            12'd 860: y = 16'hFFFF;
            12'd 861: y = 16'hFFFF;
            12'd 862: y = 16'hFFFF;
            12'd 863: y = 16'hFFFF;
            12'd 864: y = 16'hFFFF;
            12'd 865: y = 16'hFFFF;
            12'd 866: y = 16'hFFFF;
            12'd 867: y = 16'hFFFF;
            12'd 868: y = 16'hFFFF;
            12'd 869: y = 16'hFFFF;
            12'd 870: y = 16'hFFFF;
            12'd 871: y = 16'hFFFF;
            12'd 872: y = 16'hFFFF;
            12'd 873: y = 16'hFFFF;
            12'd 874: y = 16'hFFFF;
            12'd 875: y = 16'hFFFF;
            12'd 876: y = 16'hFFFF;
            12'd 877: y = 16'hFFFF;
            12'd 878: y = 16'hFFFF;
            12'd 879: y = 16'hFFFF;
            12'd 880: y = 16'hFFFF;
            12'd 881: y = 16'hFFFF;
            12'd 882: y = 16'hFFFF;
            12'd 883: y = 16'hFFFF;
            12'd 884: y = 16'hFFFF;
            12'd 885: y = 16'hFFFF;
            12'd 886: y = 16'hFFFF;
            12'd 887: y = 16'hFFFF;
            12'd 888: y = 16'hFFFF;
            12'd 889: y = 16'hFFFF;
            12'd 890: y = 16'hFFFF;
            12'd 891: y = 16'hFFFF;
            12'd 892: y = 16'hFFFF;
            12'd 893: y = 16'hFFFF;
            12'd 894: y = 16'hFFFF;
            12'd 895: y = 16'hFFFF;
            12'd 896: y = 16'hFFFF;
            12'd 897: y = 16'hFFFF;
            12'd 898: y = 16'hFFFF;
            12'd 899: y = 16'hFFFF;
            12'd 900: y = 16'hFFFF;
            12'd 901: y = 16'hFFFF;
            12'd 902: y = 16'hFFFF;
            12'd 903: y = 16'hFFFF;
            12'd 904: y = 16'hFFFF;
            12'd 905: y = 16'hFFFF;
            12'd 906: y = 16'hFFFF;
            12'd 907: y = 16'hFFFF;
            12'd 908: y = 16'hFFFF;
            12'd 909: y = 16'hFFFF;
            12'd 910: y = 16'hFFFF;
            12'd 911: y = 16'hFFFF;
            12'd 912: y = 16'hFFFF;
            12'd 913: y = 16'hFFFF;
            12'd 914: y = 16'hFFFF;
            12'd 915: y = 16'hFFFF;
            12'd 916: y = 16'hFFFF;
            12'd 917: y = 16'hFFFF;
            12'd 918: y = 16'hFFFF;
            12'd 919: y = 16'hFFFF;
            12'd 920: y = 16'hFFFF;
            12'd 921: y = 16'hFFFF;
            12'd 922: y = 16'hFFFF;
            12'd 923: y = 16'hFFFF;
            12'd 924: y = 16'hFFFF;
            12'd 925: y = 16'hFFFF;
            12'd 926: y = 16'hFFFF;
            12'd 927: y = 16'hFFFF;
            12'd 928: y = 16'hFFFF;
            12'd 929: y = 16'hFFFF;
            12'd 930: y = 16'hFFFF;
            12'd 931: y = 16'hFFFF;
            12'd 932: y = 16'hFFFF;
            12'd 933: y = 16'hFFFF;
            12'd 934: y = 16'hFFFF;
            12'd 935: y = 16'hFFFF;
            12'd 936: y = 16'hFFFF;
            12'd 937: y = 16'hFFFF;
            12'd 938: y = 16'hFFFF;
            12'd 939: y = 16'hFFFF;
            12'd 940: y = 16'hFFFF;
            12'd 941: y = 16'hFFFF;
            12'd 942: y = 16'hFFFF;
            12'd 943: y = 16'hFFFF;
            12'd 944: y = 16'hFFFF;
            12'd 945: y = 16'hFFFF;
            12'd 946: y = 16'hFFFF;
            12'd 947: y = 16'hFFFF;
            12'd 948: y = 16'hFFFF;
            12'd 949: y = 16'hFFFF;
            12'd 950: y = 16'hFFFF;
            12'd 951: y = 16'hFFFF;
            12'd 952: y = 16'hFFFF;
            12'd 953: y = 16'hFFFF;
            12'd 954: y = 16'hFFFF;
            12'd 955: y = 16'hFFFF;
            12'd 956: y = 16'hFFFF;
            12'd 957: y = 16'hFFFF;
            12'd 958: y = 16'hFFFF;
            12'd 959: y = 16'hFFFF;
            12'd 960: y = 16'hFFFF;
            12'd 961: y = 16'hFFFF;
            12'd 962: y = 16'hFFFF;
            12'd 963: y = 16'hFFFF;
            12'd 964: y = 16'hFFFF;
            12'd 965: y = 16'hFFFF;
            12'd 966: y = 16'hFFFF;
            12'd 967: y = 16'hFFFF;
            12'd 968: y = 16'hFFFF;
            12'd 969: y = 16'hFFFF;
            12'd 970: y = 16'hFFFF;
            12'd 971: y = 16'hFFFF;
            12'd 972: y = 16'hFFFF;
            12'd 973: y = 16'hFFFF;
            12'd 974: y = 16'hFFFF;
            12'd 975: y = 16'hFFFF;
            12'd 976: y = 16'hFFFF;
            12'd 977: y = 16'hFFFF;
            12'd 978: y = 16'hFFFF;
            12'd 979: y = 16'hFFFF;
            12'd 980: y = 16'hFFFF;
            12'd 981: y = 16'hFFFF;
            12'd 982: y = 16'hFFFF;
            12'd 983: y = 16'hFFFF;
            12'd 984: y = 16'hFFFF;
            12'd 985: y = 16'hFFFF;
            12'd 986: y = 16'hFFFF;
            12'd 987: y = 16'hFFFF;
            12'd 988: y = 16'hFFFF;
            12'd 989: y = 16'hFFFF;
            12'd 990: y = 16'hFFFF;
            12'd 991: y = 16'hFFFF;
            12'd 992: y = 16'hFFFF;
            12'd 993: y = 16'hFFFF;
            12'd 994: y = 16'hFFFF;
            12'd 995: y = 16'hFFFF;
            12'd 996: y = 16'hFFFF;
            12'd 997: y = 16'hFFFF;
            12'd 998: y = 16'hFFFF;
            12'd 999: y = 16'hFFFF;
            12'd1000: y = 16'hFFFF;
            12'd1001: y = 16'hFFFF;
            12'd1002: y = 16'hFFFF;
            12'd1003: y = 16'hFFFF;
            12'd1004: y = 16'hFFFF;
            12'd1005: y = 16'hFFFF;
            12'd1006: y = 16'hFFFF;
            12'd1007: y = 16'hFFFF;
            12'd1008: y = 16'hFFFF;
            12'd1009: y = 16'hFFFF;
            12'd1010: y = 16'hFFFF;
            12'd1011: y = 16'hFFFF;
            12'd1012: y = 16'hFFFF;
            12'd1013: y = 16'hFFFF;
            12'd1014: y = 16'hFFFF;
            12'd1015: y = 16'hFFFF;
            12'd1016: y = 16'hFFFF;
            12'd1017: y = 16'hFFFF;
            12'd1018: y = 16'hFFFF;
            12'd1019: y = 16'hFFFF;
            12'd1020: y = 16'hFFFF;
            12'd1021: y = 16'hFFFF;
            12'd1022: y = 16'hFFFF;
            12'd1023: y = 16'hFFFF;
            12'd1024: y = 16'hFFFF;
            12'd1025: y = 16'hFFC0;
            12'd1026: y = 16'hFF80;
            12'd1027: y = 16'hFF41;
            12'd1028: y = 16'hFF01;
            12'd1029: y = 16'hFEC2;
            12'd1030: y = 16'hFE82;
            12'd1031: y = 16'hFE43;
            12'd1032: y = 16'hFE04;
            12'd1033: y = 16'hFDC5;
            12'd1034: y = 16'hFD86;
            12'd1035: y = 16'hFD47;
            12'd1036: y = 16'hFD09;
            12'd1037: y = 16'hFCCA;
            12'd1038: y = 16'hFC8C;
            12'd1039: y = 16'hFC4E;
            12'd1040: y = 16'hFC10;
            12'd1041: y = 16'hFBD2;
            12'd1042: y = 16'hFB94;
            12'd1043: y = 16'hFB56;
            12'd1044: y = 16'hFB19;
            12'd1045: y = 16'hFADB;
            12'd1046: y = 16'hFA9E;
            12'd1047: y = 16'hFA60;
            12'd1048: y = 16'hFA23;
            12'd1049: y = 16'hF9E6;
            12'd1050: y = 16'hF9A9;
            12'd1051: y = 16'hF96C;
            12'd1052: y = 16'hF930;
            12'd1053: y = 16'hF8F3;
            12'd1054: y = 16'hF8B7;
            12'd1055: y = 16'hF87A;
            12'd1056: y = 16'hF83E;
            12'd1057: y = 16'hF802;
            12'd1058: y = 16'hF7C6;
            12'd1059: y = 16'hF78A;
            12'd1060: y = 16'hF74E;
            12'd1061: y = 16'hF713;
            12'd1062: y = 16'hF6D7;
            12'd1063: y = 16'hF69C;
            12'd1064: y = 16'hF660;
            12'd1065: y = 16'hF625;
            12'd1066: y = 16'hF5EA;
            12'd1067: y = 16'hF5AF;
            12'd1068: y = 16'hF574;
            12'd1069: y = 16'hF539;
            12'd1070: y = 16'hF4FF;
            12'd1071: y = 16'hF4C4;
            12'd1072: y = 16'hF48A;
            12'd1073: y = 16'hF44F;
            12'd1074: y = 16'hF415;
            12'd1075: y = 16'hF3DB;
            12'd1076: y = 16'hF3A1;
            12'd1077: y = 16'hF367;
            12'd1078: y = 16'hF32D;
            12'd1079: y = 16'hF2F3;
            12'd1080: y = 16'hF2BA;
            12'd1081: y = 16'hF280;
            12'd1082: y = 16'hF247;
            12'd1083: y = 16'hF20E;
            12'd1084: y = 16'hF1D5;
            12'd1085: y = 16'hF19B;
            12'd1086: y = 16'hF163;
            12'd1087: y = 16'hF12A;
            12'd1088: y = 16'hF0F1;
            12'd1089: y = 16'hF0B8;
            12'd1090: y = 16'hF080;
            12'd1091: y = 16'hF047;
            12'd1092: y = 16'hF00F;
            12'd1093: y = 16'hEFD7;
            12'd1094: y = 16'hEF9F;
            12'd1095: y = 16'hEF67;
            12'd1096: y = 16'hEF2F;
            12'd1097: y = 16'hEEF7;
            12'd1098: y = 16'hEEBF;
            12'd1099: y = 16'hEE88;
            12'd1100: y = 16'hEE50;
            12'd1101: y = 16'hEE19;
            12'd1102: y = 16'hEDE1;
            12'd1103: y = 16'hEDAA;
            12'd1104: y = 16'hED73;
            12'd1105: y = 16'hED3C;
            12'd1106: y = 16'hED05;
            12'd1107: y = 16'hECCE;
            12'd1108: y = 16'hEC98;
            12'd1109: y = 16'hEC61;
            12'd1110: y = 16'hEC2A;
            12'd1111: y = 16'hEBF4;
            12'd1112: y = 16'hEBBE;
            12'd1113: y = 16'hEB87;
            12'd1114: y = 16'hEB51;
            12'd1115: y = 16'hEB1B;
            12'd1116: y = 16'hEAE5;
            12'd1117: y = 16'hEAB0;
            12'd1118: y = 16'hEA7A;
            12'd1119: y = 16'hEA44;
            12'd1120: y = 16'hEA0F;
            12'd1121: y = 16'hE9D9;
            12'd1122: y = 16'hE9A4;
            12'd1123: y = 16'hE96F;
            12'd1124: y = 16'hE939;
            12'd1125: y = 16'hE904;
            12'd1126: y = 16'hE8CF;
            12'd1127: y = 16'hE89A;
            12'd1128: y = 16'hE866;
            12'd1129: y = 16'hE831;
            12'd1130: y = 16'hE7FC;
            12'd1131: y = 16'hE7C8;
            12'd1132: y = 16'hE793;
            12'd1133: y = 16'hE75F;
            12'd1134: y = 16'hE72B;
            12'd1135: y = 16'hE6F7;
            12'd1136: y = 16'hE6C3;
            12'd1137: y = 16'hE68F;
            12'd1138: y = 16'hE65B;
            12'd1139: y = 16'hE627;
            12'd1140: y = 16'hE5F3;
            12'd1141: y = 16'hE5C0;
            12'd1142: y = 16'hE58C;
            12'd1143: y = 16'hE559;
            12'd1144: y = 16'hE526;
            12'd1145: y = 16'hE4F2;
            12'd1146: y = 16'hE4BF;
            12'd1147: y = 16'hE48C;
            12'd1148: y = 16'hE459;
            12'd1149: y = 16'hE426;
            12'd1150: y = 16'hE3F4;
            12'd1151: y = 16'hE3C1;
            12'd1152: y = 16'hE38E;
            12'd1153: y = 16'hE35C;
            12'd1154: y = 16'hE329;
            12'd1155: y = 16'hE2F7;
            12'd1156: y = 16'hE2C5;
            12'd1157: y = 16'hE292;
            12'd1158: y = 16'hE260;
            12'd1159: y = 16'hE22E;
            12'd1160: y = 16'hE1FC;
            12'd1161: y = 16'hE1CB;
            12'd1162: y = 16'hE199;
            12'd1163: y = 16'hE167;
            12'd1164: y = 16'hE136;
            12'd1165: y = 16'hE104;
            12'd1166: y = 16'hE0D3;
            12'd1167: y = 16'hE0A1;
            12'd1168: y = 16'hE070;
            12'd1169: y = 16'hE03F;
            12'd1170: y = 16'hE00E;
            12'd1171: y = 16'hDFDD;
            12'd1172: y = 16'hDFAC;
            12'd1173: y = 16'hDF7B;
            12'd1174: y = 16'hDF4B;
            12'd1175: y = 16'hDF1A;
            12'd1176: y = 16'hDEE9;
            12'd1177: y = 16'hDEB9;
            12'd1178: y = 16'hDE88;
            12'd1179: y = 16'hDE58;
            12'd1180: y = 16'hDE28;
            12'd1181: y = 16'hDDF8;
            12'd1182: y = 16'hDDC8;
            12'd1183: y = 16'hDD98;
            12'd1184: y = 16'hDD68;
            12'd1185: y = 16'hDD38;
            12'd1186: y = 16'hDD08;
            12'd1187: y = 16'hDCD9;
            12'd1188: y = 16'hDCA9;
            12'd1189: y = 16'hDC79;
            12'd1190: y = 16'hDC4A;
            12'd1191: y = 16'hDC1B;
            12'd1192: y = 16'hDBEB;
            12'd1193: y = 16'hDBBC;
            12'd1194: y = 16'hDB8D;
            12'd1195: y = 16'hDB5E;
            12'd1196: y = 16'hDB2F;
            12'd1197: y = 16'hDB00;
            12'd1198: y = 16'hDAD1;
            12'd1199: y = 16'hDAA3;
            12'd1200: y = 16'hDA74;
            12'd1201: y = 16'hDA45;
            12'd1202: y = 16'hDA17;
            12'd1203: y = 16'hD9E9;
            12'd1204: y = 16'hD9BA;
            12'd1205: y = 16'hD98C;
            12'd1206: y = 16'hD95E;
            12'd1207: y = 16'hD930;
            12'd1208: y = 16'hD902;
            12'd1209: y = 16'hD8D4;
            12'd1210: y = 16'hD8A6;
            12'd1211: y = 16'hD878;
            12'd1212: y = 16'hD84A;
            12'd1213: y = 16'hD81D;
            12'd1214: y = 16'hD7EF;
            12'd1215: y = 16'hD7C2;
            12'd1216: y = 16'hD794;
            12'd1217: y = 16'hD767;
            12'd1218: y = 16'hD73A;
            12'd1219: y = 16'hD70C;
            12'd1220: y = 16'hD6DF;
            12'd1221: y = 16'hD6B2;
            12'd1222: y = 16'hD685;
            12'd1223: y = 16'hD658;
            12'd1224: y = 16'hD62C;
            12'd1225: y = 16'hD5FF;
            12'd1226: y = 16'hD5D2;
            12'd1227: y = 16'hD5A5;
            12'd1228: y = 16'hD579;
            12'd1229: y = 16'hD54C;
            12'd1230: y = 16'hD520;
            12'd1231: y = 16'hD4F4;
            12'd1232: y = 16'hD4C7;
            12'd1233: y = 16'hD49B;
            12'd1234: y = 16'hD46F;
            12'd1235: y = 16'hD443;
            12'd1236: y = 16'hD417;
            12'd1237: y = 16'hD3EB;
            12'd1238: y = 16'hD3BF;
            12'd1239: y = 16'hD394;
            12'd1240: y = 16'hD368;
            12'd1241: y = 16'hD33C;
            12'd1242: y = 16'hD311;
            12'd1243: y = 16'hD2E5;
            12'd1244: y = 16'hD2BA;
            12'd1245: y = 16'hD28F;
            12'd1246: y = 16'hD263;
            12'd1247: y = 16'hD238;
            12'd1248: y = 16'hD20D;
            12'd1249: y = 16'hD1E2;
            12'd1250: y = 16'hD1B7;
            12'd1251: y = 16'hD18C;
            12'd1252: y = 16'hD161;
            12'd1253: y = 16'hD137;
            12'd1254: y = 16'hD10C;
            12'd1255: y = 16'hD0E1;
            12'd1256: y = 16'hD0B7;
            12'd1257: y = 16'hD08C;
            12'd1258: y = 16'hD062;
            12'd1259: y = 16'hD037;
            12'd1260: y = 16'hD00D;
            12'd1261: y = 16'hCFE3;
            12'd1262: y = 16'hCFB9;
            12'd1263: y = 16'hCF8E;
            12'd1264: y = 16'hCF64;
            12'd1265: y = 16'hCF3A;
            12'd1266: y = 16'hCF11;
            12'd1267: y = 16'hCEE7;
            12'd1268: y = 16'hCEBD;
            12'd1269: y = 16'hCE93;
            12'd1270: y = 16'hCE6A;
            12'd1271: y = 16'hCE40;
            12'd1272: y = 16'hCE17;
            12'd1273: y = 16'hCDED;
            12'd1274: y = 16'hCDC4;
            12'd1275: y = 16'hCD9A;
            12'd1276: y = 16'hCD71;
            12'd1277: y = 16'hCD48;
            12'd1278: y = 16'hCD1F;
            12'd1279: y = 16'hCCF6;
            12'd1280: y = 16'hCCCD;
            12'd1281: y = 16'hCCA4;
            12'd1282: y = 16'hCC7B;
            12'd1283: y = 16'hCC52;
            12'd1284: y = 16'hCC29;
            12'd1285: y = 16'hCC01;
            12'd1286: y = 16'hCBD8;
            12'd1287: y = 16'hCBB0;
            12'd1288: y = 16'hCB87;
            12'd1289: y = 16'hCB5F;
            12'd1290: y = 16'hCB36;
            12'd1291: y = 16'hCB0E;
            12'd1292: y = 16'hCAE6;
            12'd1293: y = 16'hCABE;
            12'd1294: y = 16'hCA96;
            12'd1295: y = 16'hCA6E;
            12'd1296: y = 16'hCA46;
            12'd1297: y = 16'hCA1E;
            12'd1298: y = 16'hC9F6;
            12'd1299: y = 16'hC9CE;
            12'd1300: y = 16'hC9A6;
            12'd1301: y = 16'hC97F;
            12'd1302: y = 16'hC957;
            12'd1303: y = 16'hC92F;
            12'd1304: y = 16'hC908;
            12'd1305: y = 16'hC8E0;
            12'd1306: y = 16'hC8B9;
            12'd1307: y = 16'hC892;
            12'd1308: y = 16'hC86A;
            12'd1309: y = 16'hC843;
            12'd1310: y = 16'hC81C;
            12'd1311: y = 16'hC7F5;
            12'd1312: y = 16'hC7CE;
            12'd1313: y = 16'hC7A7;
            12'd1314: y = 16'hC780;
            12'd1315: y = 16'hC759;
            12'd1316: y = 16'hC733;
            12'd1317: y = 16'hC70C;
            12'd1318: y = 16'hC6E5;
            12'd1319: y = 16'hC6BF;
            12'd1320: y = 16'hC698;
            12'd1321: y = 16'hC672;
            12'd1322: y = 16'hC64B;
            12'd1323: y = 16'hC625;
            12'd1324: y = 16'hC5FE;
            12'd1325: y = 16'hC5D8;
            12'd1326: y = 16'hC5B2;
            12'd1327: y = 16'hC58C;
            12'd1328: y = 16'hC566;
            12'd1329: y = 16'hC540;
            12'd1330: y = 16'hC51A;
            12'd1331: y = 16'hC4F4;
            12'd1332: y = 16'hC4CE;
            12'd1333: y = 16'hC4A8;
            12'd1334: y = 16'hC482;
            12'd1335: y = 16'hC45D;
            12'd1336: y = 16'hC437;
            12'd1337: y = 16'hC412;
            12'd1338: y = 16'hC3EC;
            12'd1339: y = 16'hC3C7;
            12'd1340: y = 16'hC3A1;
            12'd1341: y = 16'hC37C;
            12'd1342: y = 16'hC357;
            12'd1343: y = 16'hC331;
            12'd1344: y = 16'hC30C;
            12'd1345: y = 16'hC2E7;
            12'd1346: y = 16'hC2C2;
            12'd1347: y = 16'hC29D;
            12'd1348: y = 16'hC278;
            12'd1349: y = 16'hC253;
            12'd1350: y = 16'hC22E;
            12'd1351: y = 16'hC209;
            12'd1352: y = 16'hC1E5;
            12'd1353: y = 16'hC1C0;
            12'd1354: y = 16'hC19B;
            12'd1355: y = 16'hC177;
            12'd1356: y = 16'hC152;
            12'd1357: y = 16'hC12E;
            12'd1358: y = 16'hC109;
            12'd1359: y = 16'hC0E5;
            12'd1360: y = 16'hC0C1;
            12'd1361: y = 16'hC09C;
            12'd1362: y = 16'hC078;
            12'd1363: y = 16'hC054;
            12'd1364: y = 16'hC030;
            12'd1365: y = 16'hC00C;
            12'd1366: y = 16'hBFE8;
            12'd1367: y = 16'hBFC4;
            12'd1368: y = 16'hBFA0;
            12'd1369: y = 16'hBF7C;
            12'd1370: y = 16'hBF59;
            12'd1371: y = 16'hBF35;
            12'd1372: y = 16'hBF11;
            12'd1373: y = 16'hBEEE;
            12'd1374: y = 16'hBECA;
            12'd1375: y = 16'hBEA6;
            12'd1376: y = 16'hBE83;
            12'd1377: y = 16'hBE60;
            12'd1378: y = 16'hBE3C;
            12'd1379: y = 16'hBE19;
            12'd1380: y = 16'hBDF6;
            12'd1381: y = 16'hBDD2;
            12'd1382: y = 16'hBDAF;
            12'd1383: y = 16'hBD8C;
            12'd1384: y = 16'hBD69;
            12'd1385: y = 16'hBD46;
            12'd1386: y = 16'hBD23;
            12'd1387: y = 16'hBD00;
            12'd1388: y = 16'hBCDD;
            12'd1389: y = 16'hBCBB;
            12'd1390: y = 16'hBC98;
            12'd1391: y = 16'hBC75;
            12'd1392: y = 16'hBC52;
            12'd1393: y = 16'hBC30;
            12'd1394: y = 16'hBC0D;
            12'd1395: y = 16'hBBEB;
            12'd1396: y = 16'hBBC8;
            12'd1397: y = 16'hBBA6;
            12'd1398: y = 16'hBB83;
            12'd1399: y = 16'hBB61;
            12'd1400: y = 16'hBB3F;
            12'd1401: y = 16'hBB1D;
            12'd1402: y = 16'hBAFB;
            12'd1403: y = 16'hBAD8;
            12'd1404: y = 16'hBAB6;
            12'd1405: y = 16'hBA94;
            12'd1406: y = 16'hBA72;
            12'd1407: y = 16'hBA50;
            12'd1408: y = 16'hBA2F;
            12'd1409: y = 16'hBA0D;
            12'd1410: y = 16'hB9EB;
            12'd1411: y = 16'hB9C9;
            12'd1412: y = 16'hB9A8;
            12'd1413: y = 16'hB986;
            12'd1414: y = 16'hB964;
            12'd1415: y = 16'hB943;
            12'd1416: y = 16'hB921;
            12'd1417: y = 16'hB900;
            12'd1418: y = 16'hB8DE;
            12'd1419: y = 16'hB8BD;
            12'd1420: y = 16'hB89C;
            12'd1421: y = 16'hB87B;
            12'd1422: y = 16'hB859;
            12'd1423: y = 16'hB838;
            12'd1424: y = 16'hB817;
            12'd1425: y = 16'hB7F6;
            12'd1426: y = 16'hB7D5;
            12'd1427: y = 16'hB7B4;
            12'd1428: y = 16'hB793;
            12'd1429: y = 16'hB772;
            12'd1430: y = 16'hB751;
            12'd1431: y = 16'hB730;
            12'd1432: y = 16'hB710;
            12'd1433: y = 16'hB6EF;
            12'd1434: y = 16'hB6CE;
            12'd1435: y = 16'hB6AE;
            12'd1436: y = 16'hB68D;
            12'd1437: y = 16'hB66D;
            12'd1438: y = 16'hB64C;
            12'd1439: y = 16'hB62C;
            12'd1440: y = 16'hB60B;
            12'd1441: y = 16'hB5EB;
            12'd1442: y = 16'hB5CB;
            12'd1443: y = 16'hB5AA;
            12'd1444: y = 16'hB58A;
            12'd1445: y = 16'hB56A;
            12'd1446: y = 16'hB54A;
            12'd1447: y = 16'hB52A;
            12'd1448: y = 16'hB50A;
            12'd1449: y = 16'hB4EA;
            12'd1450: y = 16'hB4CA;
            12'd1451: y = 16'hB4AA;
            12'd1452: y = 16'hB48A;
            12'd1453: y = 16'hB46A;
            12'd1454: y = 16'hB44B;
            12'd1455: y = 16'hB42B;
            12'd1456: y = 16'hB40B;
            12'd1457: y = 16'hB3EC;
            12'd1458: y = 16'hB3CC;
            12'd1459: y = 16'hB3AC;
            12'd1460: y = 16'hB38D;
            12'd1461: y = 16'hB36E;
            12'd1462: y = 16'hB34E;
            12'd1463: y = 16'hB32F;
            12'd1464: y = 16'hB30F;
            12'd1465: y = 16'hB2F0;
            12'd1466: y = 16'hB2D1;
            12'd1467: y = 16'hB2B2;
            12'd1468: y = 16'hB292;
            12'd1469: y = 16'hB273;
            12'd1470: y = 16'hB254;
            12'd1471: y = 16'hB235;
            12'd1472: y = 16'hB216;
            12'd1473: y = 16'hB1F7;
            12'd1474: y = 16'hB1D8;
            12'd1475: y = 16'hB1BA;
            12'd1476: y = 16'hB19B;
            12'd1477: y = 16'hB17C;
            12'd1478: y = 16'hB15D;
            12'd1479: y = 16'hB13E;
            12'd1480: y = 16'hB120;
            12'd1481: y = 16'hB101;
            12'd1482: y = 16'hB0E3;
            12'd1483: y = 16'hB0C4;
            12'd1484: y = 16'hB0A6;
            12'd1485: y = 16'hB087;
            12'd1486: y = 16'hB069;
            12'd1487: y = 16'hB04A;
            12'd1488: y = 16'hB02C;
            12'd1489: y = 16'hB00E;
            12'd1490: y = 16'hAFF0;
            12'd1491: y = 16'hAFD1;
            12'd1492: y = 16'hAFB3;
            12'd1493: y = 16'hAF95;
            12'd1494: y = 16'hAF77;
            12'd1495: y = 16'hAF59;
            12'd1496: y = 16'hAF3B;
            12'd1497: y = 16'hAF1D;
            12'd1498: y = 16'hAEFF;
            12'd1499: y = 16'hAEE1;
            12'd1500: y = 16'hAEC3;
            12'd1501: y = 16'hAEA5;
            12'd1502: y = 16'hAE88;
            12'd1503: y = 16'hAE6A;
            12'd1504: y = 16'hAE4C;
            12'd1505: y = 16'hAE2F;
            12'd1506: y = 16'hAE11;
            12'd1507: y = 16'hADF3;
            12'd1508: y = 16'hADD6;
            12'd1509: y = 16'hADB8;
            12'd1510: y = 16'hAD9B;
            12'd1511: y = 16'hAD7E;
            12'd1512: y = 16'hAD60;
            12'd1513: y = 16'hAD43;
            12'd1514: y = 16'hAD26;
            12'd1515: y = 16'hAD08;
            12'd1516: y = 16'hACEB;
            12'd1517: y = 16'hACCE;
            12'd1518: y = 16'hACB1;
            12'd1519: y = 16'hAC94;
            12'd1520: y = 16'hAC77;
            12'd1521: y = 16'hAC5A;
            12'd1522: y = 16'hAC3D;
            12'd1523: y = 16'hAC20;
            12'd1524: y = 16'hAC03;
            12'd1525: y = 16'hABE6;
            12'd1526: y = 16'hABC9;
            12'd1527: y = 16'hABAC;
            12'd1528: y = 16'hAB8F;
            12'd1529: y = 16'hAB73;
            12'd1530: y = 16'hAB56;
            12'd1531: y = 16'hAB39;
            12'd1532: y = 16'hAB1D;
            12'd1533: y = 16'hAB00;
            12'd1534: y = 16'hAAE4;
            12'd1535: y = 16'hAAC7;
            12'd1536: y = 16'hAAAB;
            12'd1537: y = 16'hAA8E;
            12'd1538: y = 16'hAA72;
            12'd1539: y = 16'hAA55;
            12'd1540: y = 16'hAA39;
            12'd1541: y = 16'hAA1D;
            12'd1542: y = 16'hAA01;
            12'd1543: y = 16'hA9E4;
            12'd1544: y = 16'hA9C8;
            12'd1545: y = 16'hA9AC;
            12'd1546: y = 16'hA990;
            12'd1547: y = 16'hA974;
            12'd1548: y = 16'hA958;
            12'd1549: y = 16'hA93C;
            12'd1550: y = 16'hA920;
            12'd1551: y = 16'hA904;
            12'd1552: y = 16'hA8E8;
            12'd1553: y = 16'hA8CC;
            12'd1554: y = 16'hA8B1;
            12'd1555: y = 16'hA895;
            12'd1556: y = 16'hA879;
            12'd1557: y = 16'hA85D;
            12'd1558: y = 16'hA842;
            12'd1559: y = 16'hA826;
            12'd1560: y = 16'hA80B;
            12'd1561: y = 16'hA7EF;
            12'd1562: y = 16'hA7D3;
            12'd1563: y = 16'hA7B8;
            12'd1564: y = 16'hA79C;
            12'd1565: y = 16'hA781;
            12'd1566: y = 16'hA766;
            12'd1567: y = 16'hA74A;
            12'd1568: y = 16'hA72F;
            12'd1569: y = 16'hA714;
            12'd1570: y = 16'hA6F8;
            12'd1571: y = 16'hA6DD;
            12'd1572: y = 16'hA6C2;
            12'd1573: y = 16'hA6A7;
            12'd1574: y = 16'hA68C;
            12'd1575: y = 16'hA671;
            12'd1576: y = 16'hA656;
            12'd1577: y = 16'hA63B;
            12'd1578: y = 16'hA620;
            12'd1579: y = 16'hA605;
            12'd1580: y = 16'hA5EA;
            12'd1581: y = 16'hA5CF;
            12'd1582: y = 16'hA5B4;
            12'd1583: y = 16'hA599;
            12'd1584: y = 16'hA57F;
            12'd1585: y = 16'hA564;
            12'd1586: y = 16'hA549;
            12'd1587: y = 16'hA52F;
            12'd1588: y = 16'hA514;
            12'd1589: y = 16'hA4F9;
            12'd1590: y = 16'hA4DF;
            12'd1591: y = 16'hA4C4;
            12'd1592: y = 16'hA4AA;
            12'd1593: y = 16'hA48F;
            12'd1594: y = 16'hA475;
            12'd1595: y = 16'hA45B;
            12'd1596: y = 16'hA440;
            12'd1597: y = 16'hA426;
            12'd1598: y = 16'hA40C;
            12'd1599: y = 16'hA3F1;
            12'd1600: y = 16'hA3D7;
            12'd1601: y = 16'hA3BD;
            12'd1602: y = 16'hA3A3;
            12'd1603: y = 16'hA389;
            12'd1604: y = 16'hA36E;
            12'd1605: y = 16'hA354;
            12'd1606: y = 16'hA33A;
            12'd1607: y = 16'hA320;
            12'd1608: y = 16'hA306;
            12'd1609: y = 16'hA2EC;
            12'd1610: y = 16'hA2D3;
            12'd1611: y = 16'hA2B9;
            12'd1612: y = 16'hA29F;
            12'd1613: y = 16'hA285;
            12'd1614: y = 16'hA26B;
            12'd1615: y = 16'hA251;
            12'd1616: y = 16'hA238;
            12'd1617: y = 16'hA21E;
            12'd1618: y = 16'hA204;
            12'd1619: y = 16'hA1EB;
            12'd1620: y = 16'hA1D1;
            12'd1621: y = 16'hA1B8;
            12'd1622: y = 16'hA19E;
            12'd1623: y = 16'hA185;
            12'd1624: y = 16'hA16B;
            12'd1625: y = 16'hA152;
            12'd1626: y = 16'hA138;
            12'd1627: y = 16'hA11F;
            12'd1628: y = 16'hA106;
            12'd1629: y = 16'hA0EC;
            12'd1630: y = 16'hA0D3;
            12'd1631: y = 16'hA0BA;
            12'd1632: y = 16'hA0A1;
            12'd1633: y = 16'hA087;
            12'd1634: y = 16'hA06E;
            12'd1635: y = 16'hA055;
            12'd1636: y = 16'hA03C;
            12'd1637: y = 16'hA023;
            12'd1638: y = 16'hA00A;
            12'd1639: y = 16'h9FF1;
            12'd1640: y = 16'h9FD8;
            12'd1641: y = 16'h9FBF;
            12'd1642: y = 16'h9FA6;
            12'd1643: y = 16'h9F8D;
            12'd1644: y = 16'h9F74;
            12'd1645: y = 16'h9F5C;
            12'd1646: y = 16'h9F43;
            12'd1647: y = 16'h9F2A;
            12'd1648: y = 16'h9F11;
            12'd1649: y = 16'h9EF9;
            12'd1650: y = 16'h9EE0;
            12'd1651: y = 16'h9EC7;
            12'd1652: y = 16'h9EAF;
            12'd1653: y = 16'h9E96;
            12'd1654: y = 16'h9E7E;
            12'd1655: y = 16'h9E65;
            12'd1656: y = 16'h9E4D;
            12'd1657: y = 16'h9E34;
            12'd1658: y = 16'h9E1C;
            12'd1659: y = 16'h9E03;
            12'd1660: y = 16'h9DEB;
            12'd1661: y = 16'h9DD3;
            12'd1662: y = 16'h9DBA;
            12'd1663: y = 16'h9DA2;
            12'd1664: y = 16'h9D8A;
            12'd1665: y = 16'h9D72;
            12'd1666: y = 16'h9D59;
            12'd1667: y = 16'h9D41;
            12'd1668: y = 16'h9D29;
            12'd1669: y = 16'h9D11;
            12'd1670: y = 16'h9CF9;
            12'd1671: y = 16'h9CE1;
            12'd1672: y = 16'h9CC9;
            12'd1673: y = 16'h9CB1;
            12'd1674: y = 16'h9C99;
            12'd1675: y = 16'h9C81;
            12'd1676: y = 16'h9C69;
            12'd1677: y = 16'h9C51;
            12'd1678: y = 16'h9C39;
            12'd1679: y = 16'h9C22;
            12'd1680: y = 16'h9C0A;
            12'd1681: y = 16'h9BF2;
            12'd1682: y = 16'h9BDA;
            12'd1683: y = 16'h9BC3;
            12'd1684: y = 16'h9BAB;
            12'd1685: y = 16'h9B93;
            12'd1686: y = 16'h9B7C;
            12'd1687: y = 16'h9B64;
            12'd1688: y = 16'h9B4C;
            12'd1689: y = 16'h9B35;
            12'd1690: y = 16'h9B1D;
            12'd1691: y = 16'h9B06;
            12'd1692: y = 16'h9AEE;
            12'd1693: y = 16'h9AD7;
            12'd1694: y = 16'h9AC0;
            12'd1695: y = 16'h9AA8;
            12'd1696: y = 16'h9A91;
            12'd1697: y = 16'h9A7A;
            12'd1698: y = 16'h9A62;
            12'd1699: y = 16'h9A4B;
            12'd1700: y = 16'h9A34;
            12'd1701: y = 16'h9A1D;
            12'd1702: y = 16'h9A05;
            12'd1703: y = 16'h99EE;
            12'd1704: y = 16'h99D7;
            12'd1705: y = 16'h99C0;
            12'd1706: y = 16'h99A9;
            12'd1707: y = 16'h9992;
            12'd1708: y = 16'h997B;
            12'd1709: y = 16'h9964;
            12'd1710: y = 16'h994D;
            12'd1711: y = 16'h9936;
            12'd1712: y = 16'h991F;
            12'd1713: y = 16'h9908;
            12'd1714: y = 16'h98F1;
            12'd1715: y = 16'h98DB;
            12'd1716: y = 16'h98C4;
            12'd1717: y = 16'h98AD;
            12'd1718: y = 16'h9896;
            12'd1719: y = 16'h987F;
            12'd1720: y = 16'h9869;
            12'd1721: y = 16'h9852;
            12'd1722: y = 16'h983B;
            12'd1723: y = 16'h9825;
            12'd1724: y = 16'h980E;
            12'd1725: y = 16'h97F8;
            12'd1726: y = 16'h97E1;
            12'd1727: y = 16'h97CB;
            12'd1728: y = 16'h97B4;
            12'd1729: y = 16'h979E;
            12'd1730: y = 16'h9787;
            12'd1731: y = 16'h9771;
            12'd1732: y = 16'h975A;
            12'd1733: y = 16'h9744;
            12'd1734: y = 16'h972E;
            12'd1735: y = 16'h9717;
            12'd1736: y = 16'h9701;
            12'd1737: y = 16'h96EB;
            12'd1738: y = 16'h96D5;
            12'd1739: y = 16'h96BE;
            12'd1740: y = 16'h96A8;
            12'd1741: y = 16'h9692;
            12'd1742: y = 16'h967C;
            12'd1743: y = 16'h9666;
            12'd1744: y = 16'h9650;
            12'd1745: y = 16'h963A;
            12'd1746: y = 16'h9624;
            12'd1747: y = 16'h960E;
            12'd1748: y = 16'h95F8;
            12'd1749: y = 16'h95E2;
            12'd1750: y = 16'h95CC;
            12'd1751: y = 16'h95B6;
            12'd1752: y = 16'h95A0;
            12'd1753: y = 16'h958A;
            12'd1754: y = 16'h9574;
            12'd1755: y = 16'h955F;
            12'd1756: y = 16'h9549;
            12'd1757: y = 16'h9533;
            12'd1758: y = 16'h951D;
            12'd1759: y = 16'h9508;
            12'd1760: y = 16'h94F2;
            12'd1761: y = 16'h94DC;
            12'd1762: y = 16'h94C7;
            12'd1763: y = 16'h94B1;
            12'd1764: y = 16'h949C;
            12'd1765: y = 16'h9486;
            12'd1766: y = 16'h9470;
            12'd1767: y = 16'h945B;
            12'd1768: y = 16'h9446;
            12'd1769: y = 16'h9430;
            12'd1770: y = 16'h941B;
            12'd1771: y = 16'h9405;
            12'd1772: y = 16'h93F0;
            12'd1773: y = 16'h93DA;
            12'd1774: y = 16'h93C5;
            12'd1775: y = 16'h93B0;
            12'd1776: y = 16'h939B;
            12'd1777: y = 16'h9385;
            12'd1778: y = 16'h9370;
            12'd1779: y = 16'h935B;
            12'd1780: y = 16'h9346;
            12'd1781: y = 16'h9330;
            12'd1782: y = 16'h931B;
            12'd1783: y = 16'h9306;
            12'd1784: y = 16'h92F1;
            12'd1785: y = 16'h92DC;
            12'd1786: y = 16'h92C7;
            12'd1787: y = 16'h92B2;
            12'd1788: y = 16'h929D;
            12'd1789: y = 16'h9288;
            12'd1790: y = 16'h9273;
            12'd1791: y = 16'h925E;
            12'd1792: y = 16'h9249;
            12'd1793: y = 16'h9234;
            12'd1794: y = 16'h921F;
            12'd1795: y = 16'h920B;
            12'd1796: y = 16'h91F6;
            12'd1797: y = 16'h91E1;
            12'd1798: y = 16'h91CC;
            12'd1799: y = 16'h91B7;
            12'd1800: y = 16'h91A3;
            12'd1801: y = 16'h918E;
            12'd1802: y = 16'h9179;
            12'd1803: y = 16'h9165;
            12'd1804: y = 16'h9150;
            12'd1805: y = 16'h913B;
            12'd1806: y = 16'h9127;
            12'd1807: y = 16'h9112;
            12'd1808: y = 16'h90FE;
            12'd1809: y = 16'h90E9;
            12'd1810: y = 16'h90D5;
            12'd1811: y = 16'h90C0;
            12'd1812: y = 16'h90AC;
            12'd1813: y = 16'h9097;
            12'd1814: y = 16'h9083;
            12'd1815: y = 16'h906F;
            12'd1816: y = 16'h905A;
            12'd1817: y = 16'h9046;
            12'd1818: y = 16'h9032;
            12'd1819: y = 16'h901D;
            12'd1820: y = 16'h9009;
            12'd1821: y = 16'h8FF5;
            12'd1822: y = 16'h8FE1;
            12'd1823: y = 16'h8FCC;
            12'd1824: y = 16'h8FB8;
            12'd1825: y = 16'h8FA4;
            12'd1826: y = 16'h8F90;
            12'd1827: y = 16'h8F7C;
            12'd1828: y = 16'h8F68;
            12'd1829: y = 16'h8F54;
            12'd1830: y = 16'h8F40;
            12'd1831: y = 16'h8F2B;
            12'd1832: y = 16'h8F17;
            12'd1833: y = 16'h8F03;
            12'd1834: y = 16'h8EF0;
            12'd1835: y = 16'h8EDC;
            12'd1836: y = 16'h8EC8;
            12'd1837: y = 16'h8EB4;
            12'd1838: y = 16'h8EA0;
            12'd1839: y = 16'h8E8C;
            12'd1840: y = 16'h8E78;
            12'd1841: y = 16'h8E64;
            12'd1842: y = 16'h8E51;
            12'd1843: y = 16'h8E3D;
            12'd1844: y = 16'h8E29;
            12'd1845: y = 16'h8E15;
            12'd1846: y = 16'h8E02;
            12'd1847: y = 16'h8DEE;
            12'd1848: y = 16'h8DDA;
            12'd1849: y = 16'h8DC7;
            12'd1850: y = 16'h8DB3;
            12'd1851: y = 16'h8D9F;
            12'd1852: y = 16'h8D8C;
            12'd1853: y = 16'h8D78;
            12'd1854: y = 16'h8D65;
            12'd1855: y = 16'h8D51;
            12'd1856: y = 16'h8D3E;
            12'd1857: y = 16'h8D2A;
            12'd1858: y = 16'h8D17;
            12'd1859: y = 16'h8D03;
            12'd1860: y = 16'h8CF0;
            12'd1861: y = 16'h8CDD;
            12'd1862: y = 16'h8CC9;
            12'd1863: y = 16'h8CB6;
            12'd1864: y = 16'h8CA3;
            12'd1865: y = 16'h8C8F;
            12'd1866: y = 16'h8C7C;
            12'd1867: y = 16'h8C69;
            12'd1868: y = 16'h8C56;
            12'd1869: y = 16'h8C42;
            12'd1870: y = 16'h8C2F;
            12'd1871: y = 16'h8C1C;
            12'd1872: y = 16'h8C09;
            12'd1873: y = 16'h8BF6;
            12'd1874: y = 16'h8BE2;
            12'd1875: y = 16'h8BCF;
            12'd1876: y = 16'h8BBC;
            12'd1877: y = 16'h8BA9;
            12'd1878: y = 16'h8B96;
            12'd1879: y = 16'h8B83;
            12'd1880: y = 16'h8B70;
            12'd1881: y = 16'h8B5D;
            12'd1882: y = 16'h8B4A;
            12'd1883: y = 16'h8B37;
            12'd1884: y = 16'h8B24;
            12'd1885: y = 16'h8B12;
            12'd1886: y = 16'h8AFF;
            12'd1887: y = 16'h8AEC;
            12'd1888: y = 16'h8AD9;
            12'd1889: y = 16'h8AC6;
            12'd1890: y = 16'h8AB3;
            12'd1891: y = 16'h8AA1;
            12'd1892: y = 16'h8A8E;
            12'd1893: y = 16'h8A7B;
            12'd1894: y = 16'h8A68;
            12'd1895: y = 16'h8A56;
            12'd1896: y = 16'h8A43;
            12'd1897: y = 16'h8A30;
            12'd1898: y = 16'h8A1E;
            12'd1899: y = 16'h8A0B;
            12'd1900: y = 16'h89F8;
            12'd1901: y = 16'h89E6;
            12'd1902: y = 16'h89D3;
            12'd1903: y = 16'h89C1;
            12'd1904: y = 16'h89AE;
            12'd1905: y = 16'h899C;
            12'd1906: y = 16'h8989;
            12'd1907: y = 16'h8977;
            12'd1908: y = 16'h8964;
            12'd1909: y = 16'h8952;
            12'd1910: y = 16'h8940;
            12'd1911: y = 16'h892D;
            12'd1912: y = 16'h891B;
            12'd1913: y = 16'h8908;
            12'd1914: y = 16'h88F6;
            12'd1915: y = 16'h88E4;
            12'd1916: y = 16'h88D2;
            12'd1917: y = 16'h88BF;
            12'd1918: y = 16'h88AD;
            12'd1919: y = 16'h889B;
            12'd1920: y = 16'h8889;
            12'd1921: y = 16'h8876;
            12'd1922: y = 16'h8864;
            12'd1923: y = 16'h8852;
            12'd1924: y = 16'h8840;
            12'd1925: y = 16'h882E;
            12'd1926: y = 16'h881C;
            12'd1927: y = 16'h880A;
            12'd1928: y = 16'h87F8;
            12'd1929: y = 16'h87E5;
            12'd1930: y = 16'h87D3;
            12'd1931: y = 16'h87C1;
            12'd1932: y = 16'h87AF;
            12'd1933: y = 16'h879D;
            12'd1934: y = 16'h878C;
            12'd1935: y = 16'h877A;
            12'd1936: y = 16'h8768;
            12'd1937: y = 16'h8756;
            12'd1938: y = 16'h8744;
            12'd1939: y = 16'h8732;
            12'd1940: y = 16'h8720;
            12'd1941: y = 16'h870E;
            12'd1942: y = 16'h86FD;
            12'd1943: y = 16'h86EB;
            12'd1944: y = 16'h86D9;
            12'd1945: y = 16'h86C7;
            12'd1946: y = 16'h86B6;
            12'd1947: y = 16'h86A4;
            12'd1948: y = 16'h8692;
            12'd1949: y = 16'h8680;
            12'd1950: y = 16'h866F;
            12'd1951: y = 16'h865D;
            12'd1952: y = 16'h864C;
            12'd1953: y = 16'h863A;
            12'd1954: y = 16'h8628;
            12'd1955: y = 16'h8617;
            12'd1956: y = 16'h8605;
            12'd1957: y = 16'h85F4;
            12'd1958: y = 16'h85E2;
            12'd1959: y = 16'h85D1;
            12'd1960: y = 16'h85BF;
            12'd1961: y = 16'h85AE;
            12'd1962: y = 16'h859C;
            12'd1963: y = 16'h858B;
            12'd1964: y = 16'h8579;
            12'd1965: y = 16'h8568;
            12'd1966: y = 16'h8557;
            12'd1967: y = 16'h8545;
            12'd1968: y = 16'h8534;
            12'd1969: y = 16'h8523;
            12'd1970: y = 16'h8511;
            12'd1971: y = 16'h8500;
            12'd1972: y = 16'h84EF;
            12'd1973: y = 16'h84DE;
            12'd1974: y = 16'h84CC;
            12'd1975: y = 16'h84BB;
            12'd1976: y = 16'h84AA;
            12'd1977: y = 16'h8499;
            12'd1978: y = 16'h8488;
            12'd1979: y = 16'h8476;
            12'd1980: y = 16'h8465;
            12'd1981: y = 16'h8454;
            12'd1982: y = 16'h8443;
            12'd1983: y = 16'h8432;
            12'd1984: y = 16'h8421;
            12'd1985: y = 16'h8410;
            12'd1986: y = 16'h83FF;
            12'd1987: y = 16'h83EE;
            12'd1988: y = 16'h83DD;
            12'd1989: y = 16'h83CC;
            12'd1990: y = 16'h83BB;
            12'd1991: y = 16'h83AA;
            12'd1992: y = 16'h8399;
            12'd1993: y = 16'h8388;
            12'd1994: y = 16'h8377;
            12'd1995: y = 16'h8367;
            12'd1996: y = 16'h8356;
            12'd1997: y = 16'h8345;
            12'd1998: y = 16'h8334;
            12'd1999: y = 16'h8323;
            12'd2000: y = 16'h8312;
            12'd2001: y = 16'h8302;
            12'd2002: y = 16'h82F1;
            12'd2003: y = 16'h82E0;
            12'd2004: y = 16'h82CF;
            12'd2005: y = 16'h82BF;
            12'd2006: y = 16'h82AE;
            12'd2007: y = 16'h829D;
            12'd2008: y = 16'h828D;
            12'd2009: y = 16'h827C;
            12'd2010: y = 16'h826B;
            12'd2011: y = 16'h825B;
            12'd2012: y = 16'h824A;
            12'd2013: y = 16'h823A;
            12'd2014: y = 16'h8229;
            12'd2015: y = 16'h8219;
            12'd2016: y = 16'h8208;
            12'd2017: y = 16'h81F8;
            12'd2018: y = 16'h81E7;
            12'd2019: y = 16'h81D7;
            12'd2020: y = 16'h81C6;
            12'd2021: y = 16'h81B6;
            12'd2022: y = 16'h81A5;
            12'd2023: y = 16'h8195;
            12'd2024: y = 16'h8185;
            12'd2025: y = 16'h8174;
            12'd2026: y = 16'h8164;
            12'd2027: y = 16'h8153;
            12'd2028: y = 16'h8143;
            12'd2029: y = 16'h8133;
            12'd2030: y = 16'h8123;
            12'd2031: y = 16'h8112;
            12'd2032: y = 16'h8102;
            12'd2033: y = 16'h80F2;
            12'd2034: y = 16'h80E2;
            12'd2035: y = 16'h80D1;
            12'd2036: y = 16'h80C1;
            12'd2037: y = 16'h80B1;
            12'd2038: y = 16'h80A1;
            12'd2039: y = 16'h8091;
            12'd2040: y = 16'h8081;
            12'd2041: y = 16'h8070;
            12'd2042: y = 16'h8060;
            12'd2043: y = 16'h8050;
            12'd2044: y = 16'h8040;
            12'd2045: y = 16'h8030;
            12'd2046: y = 16'h8020;
            12'd2047: y = 16'h8010;
            12'd2048: y = 16'h8000;
            12'd2049: y = 16'h7FF0;
            12'd2050: y = 16'h7FE0;
            12'd2051: y = 16'h7FD0;
            12'd2052: y = 16'h7FC0;
            12'd2053: y = 16'h7FB0;
            12'd2054: y = 16'h7FA0;
            12'd2055: y = 16'h7F90;
            12'd2056: y = 16'h7F80;
            12'd2057: y = 16'h7F71;
            12'd2058: y = 16'h7F61;
            12'd2059: y = 16'h7F51;
            12'd2060: y = 16'h7F41;
            12'd2061: y = 16'h7F31;
            12'd2062: y = 16'h7F22;
            12'd2063: y = 16'h7F12;
            12'd2064: y = 16'h7F02;
            12'd2065: y = 16'h7EF2;
            12'd2066: y = 16'h7EE3;
            12'd2067: y = 16'h7ED3;
            12'd2068: y = 16'h7EC3;
            12'd2069: y = 16'h7EB3;
            12'd2070: y = 16'h7EA4;
            12'd2071: y = 16'h7E94;
            12'd2072: y = 16'h7E84;
            12'd2073: y = 16'h7E75;
            12'd2074: y = 16'h7E65;
            12'd2075: y = 16'h7E56;
            12'd2076: y = 16'h7E46;
            12'd2077: y = 16'h7E36;
            12'd2078: y = 16'h7E27;
            12'd2079: y = 16'h7E17;
            12'd2080: y = 16'h7E08;
            12'd2081: y = 16'h7DF8;
            12'd2082: y = 16'h7DE9;
            12'd2083: y = 16'h7DD9;
            12'd2084: y = 16'h7DCA;
            12'd2085: y = 16'h7DBB;
            12'd2086: y = 16'h7DAB;
            12'd2087: y = 16'h7D9C;
            12'd2088: y = 16'h7D8C;
            12'd2089: y = 16'h7D7D;
            12'd2090: y = 16'h7D6E;
            12'd2091: y = 16'h7D5E;
            12'd2092: y = 16'h7D4F;
            12'd2093: y = 16'h7D3F;
            12'd2094: y = 16'h7D30;
            12'd2095: y = 16'h7D21;
            12'd2096: y = 16'h7D12;
            12'd2097: y = 16'h7D02;
            12'd2098: y = 16'h7CF3;
            12'd2099: y = 16'h7CE4;
            12'd2100: y = 16'h7CD5;
            12'd2101: y = 16'h7CC5;
            12'd2102: y = 16'h7CB6;
            12'd2103: y = 16'h7CA7;
            12'd2104: y = 16'h7C98;
            12'd2105: y = 16'h7C89;
            12'd2106: y = 16'h7C7A;
            12'd2107: y = 16'h7C6A;
            12'd2108: y = 16'h7C5B;
            12'd2109: y = 16'h7C4C;
            12'd2110: y = 16'h7C3D;
            12'd2111: y = 16'h7C2E;
            12'd2112: y = 16'h7C1F;
            12'd2113: y = 16'h7C10;
            12'd2114: y = 16'h7C01;
            12'd2115: y = 16'h7BF2;
            12'd2116: y = 16'h7BE3;
            12'd2117: y = 16'h7BD4;
            12'd2118: y = 16'h7BC5;
            12'd2119: y = 16'h7BB6;
            12'd2120: y = 16'h7BA7;
            12'd2121: y = 16'h7B98;
            12'd2122: y = 16'h7B89;
            12'd2123: y = 16'h7B7A;
            12'd2124: y = 16'h7B6C;
            12'd2125: y = 16'h7B5D;
            12'd2126: y = 16'h7B4E;
            12'd2127: y = 16'h7B3F;
            12'd2128: y = 16'h7B30;
            12'd2129: y = 16'h7B21;
            12'd2130: y = 16'h7B13;
            12'd2131: y = 16'h7B04;
            12'd2132: y = 16'h7AF5;
            12'd2133: y = 16'h7AE6;
            12'd2134: y = 16'h7AD7;
            12'd2135: y = 16'h7AC9;
            12'd2136: y = 16'h7ABA;
            12'd2137: y = 16'h7AAB;
            12'd2138: y = 16'h7A9D;
            12'd2139: y = 16'h7A8E;
            12'd2140: y = 16'h7A7F;
            12'd2141: y = 16'h7A71;
            12'd2142: y = 16'h7A62;
            12'd2143: y = 16'h7A53;
            12'd2144: y = 16'h7A45;
            12'd2145: y = 16'h7A36;
            12'd2146: y = 16'h7A28;
            12'd2147: y = 16'h7A19;
            12'd2148: y = 16'h7A0A;
            12'd2149: y = 16'h79FC;
            12'd2150: y = 16'h79ED;
            12'd2151: y = 16'h79DF;
            12'd2152: y = 16'h79D0;
            12'd2153: y = 16'h79C2;
            12'd2154: y = 16'h79B3;
            12'd2155: y = 16'h79A5;
            12'd2156: y = 16'h7997;
            12'd2157: y = 16'h7988;
            12'd2158: y = 16'h797A;
            12'd2159: y = 16'h796B;
            12'd2160: y = 16'h795D;
            12'd2161: y = 16'h794F;
            12'd2162: y = 16'h7940;
            12'd2163: y = 16'h7932;
            12'd2164: y = 16'h7923;
            12'd2165: y = 16'h7915;
            12'd2166: y = 16'h7907;
            12'd2167: y = 16'h78F9;
            12'd2168: y = 16'h78EA;
            12'd2169: y = 16'h78DC;
            12'd2170: y = 16'h78CE;
            12'd2171: y = 16'h78BF;
            12'd2172: y = 16'h78B1;
            12'd2173: y = 16'h78A3;
            12'd2174: y = 16'h7895;
            12'd2175: y = 16'h7887;
            12'd2176: y = 16'h7878;
            12'd2177: y = 16'h786A;
            12'd2178: y = 16'h785C;
            12'd2179: y = 16'h784E;
            12'd2180: y = 16'h7840;
            12'd2181: y = 16'h7832;
            12'd2182: y = 16'h7824;
            12'd2183: y = 16'h7816;
            12'd2184: y = 16'h7808;
            12'd2185: y = 16'h77F9;
            12'd2186: y = 16'h77EB;
            12'd2187: y = 16'h77DD;
            12'd2188: y = 16'h77CF;
            12'd2189: y = 16'h77C1;
            12'd2190: y = 16'h77B3;
            12'd2191: y = 16'h77A5;
            12'd2192: y = 16'h7797;
            12'd2193: y = 16'h7789;
            12'd2194: y = 16'h777B;
            12'd2195: y = 16'h776E;
            12'd2196: y = 16'h7760;
            12'd2197: y = 16'h7752;
            12'd2198: y = 16'h7744;
            12'd2199: y = 16'h7736;
            12'd2200: y = 16'h7728;
            12'd2201: y = 16'h771A;
            12'd2202: y = 16'h770C;
            12'd2203: y = 16'h76FE;
            12'd2204: y = 16'h76F1;
            12'd2205: y = 16'h76E3;
            12'd2206: y = 16'h76D5;
            12'd2207: y = 16'h76C7;
            12'd2208: y = 16'h76BA;
            12'd2209: y = 16'h76AC;
            12'd2210: y = 16'h769E;
            12'd2211: y = 16'h7690;
            12'd2212: y = 16'h7683;
            12'd2213: y = 16'h7675;
            12'd2214: y = 16'h7667;
            12'd2215: y = 16'h7659;
            12'd2216: y = 16'h764C;
            12'd2217: y = 16'h763E;
            12'd2218: y = 16'h7630;
            12'd2219: y = 16'h7623;
            12'd2220: y = 16'h7615;
            12'd2221: y = 16'h7608;
            12'd2222: y = 16'h75FA;
            12'd2223: y = 16'h75EC;
            12'd2224: y = 16'h75DF;
            12'd2225: y = 16'h75D1;
            12'd2226: y = 16'h75C4;
            12'd2227: y = 16'h75B6;
            12'd2228: y = 16'h75A9;
            12'd2229: y = 16'h759B;
            12'd2230: y = 16'h758E;
            12'd2231: y = 16'h7580;
            12'd2232: y = 16'h7573;
            12'd2233: y = 16'h7565;
            12'd2234: y = 16'h7558;
            12'd2235: y = 16'h754A;
            12'd2236: y = 16'h753D;
            12'd2237: y = 16'h752F;
            12'd2238: y = 16'h7522;
            12'd2239: y = 16'h7515;
            12'd2240: y = 16'h7507;
            12'd2241: y = 16'h74FA;
            12'd2242: y = 16'h74ED;
            12'd2243: y = 16'h74DF;
            12'd2244: y = 16'h74D2;
            12'd2245: y = 16'h74C5;
            12'd2246: y = 16'h74B7;
            12'd2247: y = 16'h74AA;
            12'd2248: y = 16'h749D;
            12'd2249: y = 16'h748F;
            12'd2250: y = 16'h7482;
            12'd2251: y = 16'h7475;
            12'd2252: y = 16'h7468;
            12'd2253: y = 16'h745A;
            12'd2254: y = 16'h744D;
            12'd2255: y = 16'h7440;
            12'd2256: y = 16'h7433;
            12'd2257: y = 16'h7426;
            12'd2258: y = 16'h7418;
            12'd2259: y = 16'h740B;
            12'd2260: y = 16'h73FE;
            12'd2261: y = 16'h73F1;
            12'd2262: y = 16'h73E4;
            12'd2263: y = 16'h73D7;
            12'd2264: y = 16'h73CA;
            12'd2265: y = 16'h73BD;
            12'd2266: y = 16'h73B0;
            12'd2267: y = 16'h73A2;
            12'd2268: y = 16'h7395;
            12'd2269: y = 16'h7388;
            12'd2270: y = 16'h737B;
            12'd2271: y = 16'h736E;
            12'd2272: y = 16'h7361;
            12'd2273: y = 16'h7354;
            12'd2274: y = 16'h7347;
            12'd2275: y = 16'h733A;
            12'd2276: y = 16'h732D;
            12'd2277: y = 16'h7320;
            12'd2278: y = 16'h7314;
            12'd2279: y = 16'h7307;
            12'd2280: y = 16'h72FA;
            12'd2281: y = 16'h72ED;
            12'd2282: y = 16'h72E0;
            12'd2283: y = 16'h72D3;
            12'd2284: y = 16'h72C6;
            12'd2285: y = 16'h72B9;
            12'd2286: y = 16'h72AC;
            12'd2287: y = 16'h72A0;
            12'd2288: y = 16'h7293;
            12'd2289: y = 16'h7286;
            12'd2290: y = 16'h7279;
            12'd2291: y = 16'h726C;
            12'd2292: y = 16'h7260;
            12'd2293: y = 16'h7253;
            12'd2294: y = 16'h7246;
            12'd2295: y = 16'h7239;
            12'd2296: y = 16'h722D;
            12'd2297: y = 16'h7220;
            12'd2298: y = 16'h7213;
            12'd2299: y = 16'h7206;
            12'd2300: y = 16'h71FA;
            12'd2301: y = 16'h71ED;
            12'd2302: y = 16'h71E0;
            12'd2303: y = 16'h71D4;
            12'd2304: y = 16'h71C7;
            12'd2305: y = 16'h71BA;
            12'd2306: y = 16'h71AE;
            12'd2307: y = 16'h71A1;
            12'd2308: y = 16'h7195;
            12'd2309: y = 16'h7188;
            12'd2310: y = 16'h717B;
            12'd2311: y = 16'h716F;
            12'd2312: y = 16'h7162;
            12'd2313: y = 16'h7156;
            12'd2314: y = 16'h7149;
            12'd2315: y = 16'h713D;
            12'd2316: y = 16'h7130;
            12'd2317: y = 16'h7124;
            12'd2318: y = 16'h7117;
            12'd2319: y = 16'h710B;
            12'd2320: y = 16'h70FE;
            12'd2321: y = 16'h70F2;
            12'd2322: y = 16'h70E5;
            12'd2323: y = 16'h70D9;
            12'd2324: y = 16'h70CC;
            12'd2325: y = 16'h70C0;
            12'd2326: y = 16'h70B4;
            12'd2327: y = 16'h70A7;
            12'd2328: y = 16'h709B;
            12'd2329: y = 16'h708E;
            12'd2330: y = 16'h7082;
            12'd2331: y = 16'h7076;
            12'd2332: y = 16'h7069;
            12'd2333: y = 16'h705D;
            12'd2334: y = 16'h7051;
            12'd2335: y = 16'h7044;
            12'd2336: y = 16'h7038;
            12'd2337: y = 16'h702C;
            12'd2338: y = 16'h7020;
            12'd2339: y = 16'h7013;
            12'd2340: y = 16'h7007;
            12'd2341: y = 16'h6FFB;
            12'd2342: y = 16'h6FEF;
            12'd2343: y = 16'h6FE2;
            12'd2344: y = 16'h6FD6;
            12'd2345: y = 16'h6FCA;
            12'd2346: y = 16'h6FBE;
            12'd2347: y = 16'h6FB1;
            12'd2348: y = 16'h6FA5;
            12'd2349: y = 16'h6F99;
            12'd2350: y = 16'h6F8D;
            12'd2351: y = 16'h6F81;
            12'd2352: y = 16'h6F75;
            12'd2353: y = 16'h6F69;
            12'd2354: y = 16'h6F5C;
            12'd2355: y = 16'h6F50;
            12'd2356: y = 16'h6F44;
            12'd2357: y = 16'h6F38;
            12'd2358: y = 16'h6F2C;
            12'd2359: y = 16'h6F20;
            12'd2360: y = 16'h6F14;
            12'd2361: y = 16'h6F08;
            12'd2362: y = 16'h6EFC;
            12'd2363: y = 16'h6EF0;
            12'd2364: y = 16'h6EE4;
            12'd2365: y = 16'h6ED8;
            12'd2366: y = 16'h6ECC;
            12'd2367: y = 16'h6EC0;
            12'd2368: y = 16'h6EB4;
            12'd2369: y = 16'h6EA8;
            12'd2370: y = 16'h6E9C;
            12'd2371: y = 16'h6E90;
            12'd2372: y = 16'h6E84;
            12'd2373: y = 16'h6E78;
            12'd2374: y = 16'h6E6C;
            12'd2375: y = 16'h6E60;
            12'd2376: y = 16'h6E54;
            12'd2377: y = 16'h6E49;
            12'd2378: y = 16'h6E3D;
            12'd2379: y = 16'h6E31;
            12'd2380: y = 16'h6E25;
            12'd2381: y = 16'h6E19;
            12'd2382: y = 16'h6E0D;
            12'd2383: y = 16'h6E02;
            12'd2384: y = 16'h6DF6;
            12'd2385: y = 16'h6DEA;
            12'd2386: y = 16'h6DDE;
            12'd2387: y = 16'h6DD2;
            12'd2388: y = 16'h6DC7;
            12'd2389: y = 16'h6DBB;
            12'd2390: y = 16'h6DAF;
            12'd2391: y = 16'h6DA3;
            12'd2392: y = 16'h6D98;
            12'd2393: y = 16'h6D8C;
            12'd2394: y = 16'h6D80;
            12'd2395: y = 16'h6D74;
            12'd2396: y = 16'h6D69;
            12'd2397: y = 16'h6D5D;
            12'd2398: y = 16'h6D51;
            12'd2399: y = 16'h6D46;
            12'd2400: y = 16'h6D3A;
            12'd2401: y = 16'h6D2E;
            12'd2402: y = 16'h6D23;
            12'd2403: y = 16'h6D17;
            12'd2404: y = 16'h6D0C;
            12'd2405: y = 16'h6D00;
            12'd2406: y = 16'h6CF4;
            12'd2407: y = 16'h6CE9;
            12'd2408: y = 16'h6CDD;
            12'd2409: y = 16'h6CD2;
            12'd2410: y = 16'h6CC6;
            12'd2411: y = 16'h6CBA;
            12'd2412: y = 16'h6CAF;
            12'd2413: y = 16'h6CA3;
            12'd2414: y = 16'h6C98;
            12'd2415: y = 16'h6C8C;
            12'd2416: y = 16'h6C81;
            12'd2417: y = 16'h6C75;
            12'd2418: y = 16'h6C6A;
            12'd2419: y = 16'h6C5E;
            12'd2420: y = 16'h6C53;
            12'd2421: y = 16'h6C47;
            12'd2422: y = 16'h6C3C;
            12'd2423: y = 16'h6C31;
            12'd2424: y = 16'h6C25;
            12'd2425: y = 16'h6C1A;
            12'd2426: y = 16'h6C0E;
            12'd2427: y = 16'h6C03;
            12'd2428: y = 16'h6BF8;
            12'd2429: y = 16'h6BEC;
            12'd2430: y = 16'h6BE1;
            12'd2431: y = 16'h6BD5;
            12'd2432: y = 16'h6BCA;
            12'd2433: y = 16'h6BBF;
            12'd2434: y = 16'h6BB3;
            12'd2435: y = 16'h6BA8;
            12'd2436: y = 16'h6B9D;
            12'd2437: y = 16'h6B91;
            12'd2438: y = 16'h6B86;
            12'd2439: y = 16'h6B7B;
            12'd2440: y = 16'h6B70;
            12'd2441: y = 16'h6B64;
            12'd2442: y = 16'h6B59;
            12'd2443: y = 16'h6B4E;
            12'd2444: y = 16'h6B43;
            12'd2445: y = 16'h6B37;
            12'd2446: y = 16'h6B2C;
            12'd2447: y = 16'h6B21;
            12'd2448: y = 16'h6B16;
            12'd2449: y = 16'h6B0B;
            12'd2450: y = 16'h6AFF;
            12'd2451: y = 16'h6AF4;
            12'd2452: y = 16'h6AE9;
            12'd2453: y = 16'h6ADE;
            12'd2454: y = 16'h6AD3;
            12'd2455: y = 16'h6AC8;
            12'd2456: y = 16'h6ABC;
            12'd2457: y = 16'h6AB1;
            12'd2458: y = 16'h6AA6;
            12'd2459: y = 16'h6A9B;
            12'd2460: y = 16'h6A90;
            12'd2461: y = 16'h6A85;
            12'd2462: y = 16'h6A7A;
            12'd2463: y = 16'h6A6F;
            12'd2464: y = 16'h6A64;
            12'd2465: y = 16'h6A59;
            12'd2466: y = 16'h6A4E;
            12'd2467: y = 16'h6A43;
            12'd2468: y = 16'h6A38;
            12'd2469: y = 16'h6A2D;
            12'd2470: y = 16'h6A22;
            12'd2471: y = 16'h6A17;
            12'd2472: y = 16'h6A0C;
            12'd2473: y = 16'h6A01;
            12'd2474: y = 16'h69F6;
            12'd2475: y = 16'h69EB;
            12'd2476: y = 16'h69E0;
            12'd2477: y = 16'h69D5;
            12'd2478: y = 16'h69CA;
            12'd2479: y = 16'h69BF;
            12'd2480: y = 16'h69B4;
            12'd2481: y = 16'h69A9;
            12'd2482: y = 16'h699E;
            12'd2483: y = 16'h6993;
            12'd2484: y = 16'h6988;
            12'd2485: y = 16'h697E;
            12'd2486: y = 16'h6973;
            12'd2487: y = 16'h6968;
            12'd2488: y = 16'h695D;
            12'd2489: y = 16'h6952;
            12'd2490: y = 16'h6947;
            12'd2491: y = 16'h693D;
            12'd2492: y = 16'h6932;
            12'd2493: y = 16'h6927;
            12'd2494: y = 16'h691C;
            12'd2495: y = 16'h6911;
            12'd2496: y = 16'h6907;
            12'd2497: y = 16'h68FC;
            12'd2498: y = 16'h68F1;
            12'd2499: y = 16'h68E6;
            12'd2500: y = 16'h68DC;
            12'd2501: y = 16'h68D1;
            12'd2502: y = 16'h68C6;
            12'd2503: y = 16'h68BB;
            12'd2504: y = 16'h68B1;
            12'd2505: y = 16'h68A6;
            12'd2506: y = 16'h689B;
            12'd2507: y = 16'h6891;
            12'd2508: y = 16'h6886;
            12'd2509: y = 16'h687B;
            12'd2510: y = 16'h6871;
            12'd2511: y = 16'h6866;
            12'd2512: y = 16'h685B;
            12'd2513: y = 16'h6851;
            12'd2514: y = 16'h6846;
            12'd2515: y = 16'h683B;
            12'd2516: y = 16'h6831;
            12'd2517: y = 16'h6826;
            12'd2518: y = 16'h681C;
            12'd2519: y = 16'h6811;
            12'd2520: y = 16'h6807;
            12'd2521: y = 16'h67FC;
            12'd2522: y = 16'h67F1;
            12'd2523: y = 16'h67E7;
            12'd2524: y = 16'h67DC;
            12'd2525: y = 16'h67D2;
            12'd2526: y = 16'h67C7;
            12'd2527: y = 16'h67BD;
            12'd2528: y = 16'h67B2;
            12'd2529: y = 16'h67A8;
            12'd2530: y = 16'h679D;
            12'd2531: y = 16'h6793;
            12'd2532: y = 16'h6788;
            12'd2533: y = 16'h677E;
            12'd2534: y = 16'h6773;
            12'd2535: y = 16'h6769;
            12'd2536: y = 16'h675E;
            12'd2537: y = 16'h6754;
            12'd2538: y = 16'h674A;
            12'd2539: y = 16'h673F;
            12'd2540: y = 16'h6735;
            12'd2541: y = 16'h672A;
            12'd2542: y = 16'h6720;
            12'd2543: y = 16'h6716;
            12'd2544: y = 16'h670B;
            12'd2545: y = 16'h6701;
            12'd2546: y = 16'h66F7;
            12'd2547: y = 16'h66EC;
            12'd2548: y = 16'h66E2;
            12'd2549: y = 16'h66D8;
            12'd2550: y = 16'h66CD;
            12'd2551: y = 16'h66C3;
            12'd2552: y = 16'h66B9;
            12'd2553: y = 16'h66AE;
            12'd2554: y = 16'h66A4;
            12'd2555: y = 16'h669A;
            12'd2556: y = 16'h668F;
            12'd2557: y = 16'h6685;
            12'd2558: y = 16'h667B;
            12'd2559: y = 16'h6671;
            12'd2560: y = 16'h6666;
            12'd2561: y = 16'h665C;
            12'd2562: y = 16'h6652;
            12'd2563: y = 16'h6648;
            12'd2564: y = 16'h663E;
            12'd2565: y = 16'h6633;
            12'd2566: y = 16'h6629;
            12'd2567: y = 16'h661F;
            12'd2568: y = 16'h6615;
            12'd2569: y = 16'h660B;
            12'd2570: y = 16'h6600;
            12'd2571: y = 16'h65F6;
            12'd2572: y = 16'h65EC;
            12'd2573: y = 16'h65E2;
            12'd2574: y = 16'h65D8;
            12'd2575: y = 16'h65CE;
            12'd2576: y = 16'h65C4;
            12'd2577: y = 16'h65B9;
            12'd2578: y = 16'h65AF;
            12'd2579: y = 16'h65A5;
            12'd2580: y = 16'h659B;
            12'd2581: y = 16'h6591;
            12'd2582: y = 16'h6587;
            12'd2583: y = 16'h657D;
            12'd2584: y = 16'h6573;
            12'd2585: y = 16'h6569;
            12'd2586: y = 16'h655F;
            12'd2587: y = 16'h6555;
            12'd2588: y = 16'h654B;
            12'd2589: y = 16'h6541;
            12'd2590: y = 16'h6537;
            12'd2591: y = 16'h652D;
            12'd2592: y = 16'h6523;
            12'd2593: y = 16'h6519;
            12'd2594: y = 16'h650F;
            12'd2595: y = 16'h6505;
            12'd2596: y = 16'h64FB;
            12'd2597: y = 16'h64F1;
            12'd2598: y = 16'h64E7;
            12'd2599: y = 16'h64DD;
            12'd2600: y = 16'h64D3;
            12'd2601: y = 16'h64C9;
            12'd2602: y = 16'h64BF;
            12'd2603: y = 16'h64B5;
            12'd2604: y = 16'h64AB;
            12'd2605: y = 16'h64A2;
            12'd2606: y = 16'h6498;
            12'd2607: y = 16'h648E;
            12'd2608: y = 16'h6484;
            12'd2609: y = 16'h647A;
            12'd2610: y = 16'h6470;
            12'd2611: y = 16'h6466;
            12'd2612: y = 16'h645D;
            12'd2613: y = 16'h6453;
            12'd2614: y = 16'h6449;
            12'd2615: y = 16'h643F;
            12'd2616: y = 16'h6435;
            12'd2617: y = 16'h642B;
            12'd2618: y = 16'h6422;
            12'd2619: y = 16'h6418;
            12'd2620: y = 16'h640E;
            12'd2621: y = 16'h6404;
            12'd2622: y = 16'h63FB;
            12'd2623: y = 16'h63F1;
            12'd2624: y = 16'h63E7;
            12'd2625: y = 16'h63DD;
            12'd2626: y = 16'h63D4;
            12'd2627: y = 16'h63CA;
            12'd2628: y = 16'h63C0;
            12'd2629: y = 16'h63B6;
            12'd2630: y = 16'h63AD;
            12'd2631: y = 16'h63A3;
            12'd2632: y = 16'h6399;
            12'd2633: y = 16'h6390;
            12'd2634: y = 16'h6386;
            12'd2635: y = 16'h637C;
            12'd2636: y = 16'h6373;
            12'd2637: y = 16'h6369;
            12'd2638: y = 16'h635F;
            12'd2639: y = 16'h6356;
            12'd2640: y = 16'h634C;
            12'd2641: y = 16'h6342;
            12'd2642: y = 16'h6339;
            12'd2643: y = 16'h632F;
            12'd2644: y = 16'h6326;
            12'd2645: y = 16'h631C;
            12'd2646: y = 16'h6312;
            12'd2647: y = 16'h6309;
            12'd2648: y = 16'h62FF;
            12'd2649: y = 16'h62F6;
            12'd2650: y = 16'h62EC;
            12'd2651: y = 16'h62E3;
            12'd2652: y = 16'h62D9;
            12'd2653: y = 16'h62CF;
            12'd2654: y = 16'h62C6;
            12'd2655: y = 16'h62BC;
            12'd2656: y = 16'h62B3;
            12'd2657: y = 16'h62A9;
            12'd2658: y = 16'h62A0;
            12'd2659: y = 16'h6296;
            12'd2660: y = 16'h628D;
            12'd2661: y = 16'h6283;
            12'd2662: y = 16'h627A;
            12'd2663: y = 16'h6270;
            12'd2664: y = 16'h6267;
            12'd2665: y = 16'h625E;
            12'd2666: y = 16'h6254;
            12'd2667: y = 16'h624B;
            12'd2668: y = 16'h6241;
            12'd2669: y = 16'h6238;
            12'd2670: y = 16'h622E;
            12'd2671: y = 16'h6225;
            12'd2672: y = 16'h621C;
            12'd2673: y = 16'h6212;
            12'd2674: y = 16'h6209;
            12'd2675: y = 16'h61FF;
            12'd2676: y = 16'h61F6;
            12'd2677: y = 16'h61ED;
            12'd2678: y = 16'h61E3;
            12'd2679: y = 16'h61DA;
            12'd2680: y = 16'h61D1;
            12'd2681: y = 16'h61C7;
            12'd2682: y = 16'h61BE;
            12'd2683: y = 16'h61B5;
            12'd2684: y = 16'h61AB;
            12'd2685: y = 16'h61A2;
            12'd2686: y = 16'h6199;
            12'd2687: y = 16'h618F;
            12'd2688: y = 16'h6186;
            12'd2689: y = 16'h617D;
            12'd2690: y = 16'h6174;
            12'd2691: y = 16'h616A;
            12'd2692: y = 16'h6161;
            12'd2693: y = 16'h6158;
            12'd2694: y = 16'h614E;
            12'd2695: y = 16'h6145;
            12'd2696: y = 16'h613C;
            12'd2697: y = 16'h6133;
            12'd2698: y = 16'h612A;
            12'd2699: y = 16'h6120;
            12'd2700: y = 16'h6117;
            12'd2701: y = 16'h610E;
            12'd2702: y = 16'h6105;
            12'd2703: y = 16'h60FC;
            12'd2704: y = 16'h60F2;
            12'd2705: y = 16'h60E9;
            12'd2706: y = 16'h60E0;
            12'd2707: y = 16'h60D7;
            12'd2708: y = 16'h60CE;
            12'd2709: y = 16'h60C5;
            12'd2710: y = 16'h60BB;
            12'd2711: y = 16'h60B2;
            12'd2712: y = 16'h60A9;
            12'd2713: y = 16'h60A0;
            12'd2714: y = 16'h6097;
            12'd2715: y = 16'h608E;
            12'd2716: y = 16'h6085;
            12'd2717: y = 16'h607C;
            12'd2718: y = 16'h6073;
            12'd2719: y = 16'h6069;
            12'd2720: y = 16'h6060;
            12'd2721: y = 16'h6057;
            12'd2722: y = 16'h604E;
            12'd2723: y = 16'h6045;
            12'd2724: y = 16'h603C;
            12'd2725: y = 16'h6033;
            12'd2726: y = 16'h602A;
            12'd2727: y = 16'h6021;
            12'd2728: y = 16'h6018;
            12'd2729: y = 16'h600F;
            12'd2730: y = 16'h6006;
            12'd2731: y = 16'h5FFD;
            12'd2732: y = 16'h5FF4;
            12'd2733: y = 16'h5FEB;
            12'd2734: y = 16'h5FE2;
            12'd2735: y = 16'h5FD9;
            12'd2736: y = 16'h5FD0;
            12'd2737: y = 16'h5FC7;
            12'd2738: y = 16'h5FBE;
            12'd2739: y = 16'h5FB5;
            12'd2740: y = 16'h5FAC;
            12'd2741: y = 16'h5FA3;
            12'd2742: y = 16'h5F9A;
            12'd2743: y = 16'h5F91;
            12'd2744: y = 16'h5F89;
            12'd2745: y = 16'h5F80;
            12'd2746: y = 16'h5F77;
            12'd2747: y = 16'h5F6E;
            12'd2748: y = 16'h5F65;
            12'd2749: y = 16'h5F5C;
            12'd2750: y = 16'h5F53;
            12'd2751: y = 16'h5F4A;
            12'd2752: y = 16'h5F41;
            12'd2753: y = 16'h5F39;
            12'd2754: y = 16'h5F30;
            12'd2755: y = 16'h5F27;
            12'd2756: y = 16'h5F1E;
            12'd2757: y = 16'h5F15;
            12'd2758: y = 16'h5F0C;
            12'd2759: y = 16'h5F04;
            12'd2760: y = 16'h5EFB;
            12'd2761: y = 16'h5EF2;
            12'd2762: y = 16'h5EE9;
            12'd2763: y = 16'h5EE0;
            12'd2764: y = 16'h5ED8;
            12'd2765: y = 16'h5ECF;
            12'd2766: y = 16'h5EC6;
            12'd2767: y = 16'h5EBD;
            12'd2768: y = 16'h5EB5;
            12'd2769: y = 16'h5EAC;
            12'd2770: y = 16'h5EA3;
            12'd2771: y = 16'h5E9A;
            12'd2772: y = 16'h5E92;
            12'd2773: y = 16'h5E89;
            12'd2774: y = 16'h5E80;
            12'd2775: y = 16'h5E77;
            12'd2776: y = 16'h5E6F;
            12'd2777: y = 16'h5E66;
            12'd2778: y = 16'h5E5D;
            12'd2779: y = 16'h5E55;
            12'd2780: y = 16'h5E4C;
            12'd2781: y = 16'h5E43;
            12'd2782: y = 16'h5E3B;
            12'd2783: y = 16'h5E32;
            12'd2784: y = 16'h5E29;
            12'd2785: y = 16'h5E21;
            12'd2786: y = 16'h5E18;
            12'd2787: y = 16'h5E0F;
            12'd2788: y = 16'h5E07;
            12'd2789: y = 16'h5DFE;
            12'd2790: y = 16'h5DF5;
            12'd2791: y = 16'h5DED;
            12'd2792: y = 16'h5DE4;
            12'd2793: y = 16'h5DDC;
            12'd2794: y = 16'h5DD3;
            12'd2795: y = 16'h5DCA;
            12'd2796: y = 16'h5DC2;
            12'd2797: y = 16'h5DB9;
            12'd2798: y = 16'h5DB1;
            12'd2799: y = 16'h5DA8;
            12'd2800: y = 16'h5D9F;
            12'd2801: y = 16'h5D97;
            12'd2802: y = 16'h5D8E;
            12'd2803: y = 16'h5D86;
            12'd2804: y = 16'h5D7D;
            12'd2805: y = 16'h5D75;
            12'd2806: y = 16'h5D6C;
            12'd2807: y = 16'h5D64;
            12'd2808: y = 16'h5D5B;
            12'd2809: y = 16'h5D53;
            12'd2810: y = 16'h5D4A;
            12'd2811: y = 16'h5D42;
            12'd2812: y = 16'h5D39;
            12'd2813: y = 16'h5D31;
            12'd2814: y = 16'h5D28;
            12'd2815: y = 16'h5D20;
            12'd2816: y = 16'h5D17;
            12'd2817: y = 16'h5D0F;
            12'd2818: y = 16'h5D06;
            12'd2819: y = 16'h5CFE;
            12'd2820: y = 16'h5CF5;
            12'd2821: y = 16'h5CED;
            12'd2822: y = 16'h5CE5;
            12'd2823: y = 16'h5CDC;
            12'd2824: y = 16'h5CD4;
            12'd2825: y = 16'h5CCB;
            12'd2826: y = 16'h5CC3;
            12'd2827: y = 16'h5CBB;
            12'd2828: y = 16'h5CB2;
            12'd2829: y = 16'h5CAA;
            12'd2830: y = 16'h5CA1;
            12'd2831: y = 16'h5C99;
            12'd2832: y = 16'h5C91;
            12'd2833: y = 16'h5C88;
            12'd2834: y = 16'h5C80;
            12'd2835: y = 16'h5C78;
            12'd2836: y = 16'h5C6F;
            12'd2837: y = 16'h5C67;
            12'd2838: y = 16'h5C5F;
            12'd2839: y = 16'h5C56;
            12'd2840: y = 16'h5C4E;
            12'd2841: y = 16'h5C46;
            12'd2842: y = 16'h5C3D;
            12'd2843: y = 16'h5C35;
            12'd2844: y = 16'h5C2D;
            12'd2845: y = 16'h5C24;
            12'd2846: y = 16'h5C1C;
            12'd2847: y = 16'h5C14;
            12'd2848: y = 16'h5C0C;
            12'd2849: y = 16'h5C03;
            12'd2850: y = 16'h5BFB;
            12'd2851: y = 16'h5BF3;
            12'd2852: y = 16'h5BEA;
            12'd2853: y = 16'h5BE2;
            12'd2854: y = 16'h5BDA;
            12'd2855: y = 16'h5BD2;
            12'd2856: y = 16'h5BCA;
            12'd2857: y = 16'h5BC1;
            12'd2858: y = 16'h5BB9;
            12'd2859: y = 16'h5BB1;
            12'd2860: y = 16'h5BA9;
            12'd2861: y = 16'h5BA0;
            12'd2862: y = 16'h5B98;
            12'd2863: y = 16'h5B90;
            12'd2864: y = 16'h5B88;
            12'd2865: y = 16'h5B80;
            12'd2866: y = 16'h5B78;
            12'd2867: y = 16'h5B6F;
            12'd2868: y = 16'h5B67;
            12'd2869: y = 16'h5B5F;
            12'd2870: y = 16'h5B57;
            12'd2871: y = 16'h5B4F;
            12'd2872: y = 16'h5B47;
            12'd2873: y = 16'h5B3E;
            12'd2874: y = 16'h5B36;
            12'd2875: y = 16'h5B2E;
            12'd2876: y = 16'h5B26;
            12'd2877: y = 16'h5B1E;
            12'd2878: y = 16'h5B16;
            12'd2879: y = 16'h5B0E;
            12'd2880: y = 16'h5B06;
            12'd2881: y = 16'h5AFE;
            12'd2882: y = 16'h5AF6;
            12'd2883: y = 16'h5AED;
            12'd2884: y = 16'h5AE5;
            12'd2885: y = 16'h5ADD;
            12'd2886: y = 16'h5AD5;
            12'd2887: y = 16'h5ACD;
            12'd2888: y = 16'h5AC5;
            12'd2889: y = 16'h5ABD;
            12'd2890: y = 16'h5AB5;
            12'd2891: y = 16'h5AAD;
            12'd2892: y = 16'h5AA5;
            12'd2893: y = 16'h5A9D;
            12'd2894: y = 16'h5A95;
            12'd2895: y = 16'h5A8D;
            12'd2896: y = 16'h5A85;
            12'd2897: y = 16'h5A7D;
            12'd2898: y = 16'h5A75;
            12'd2899: y = 16'h5A6D;
            12'd2900: y = 16'h5A65;
            12'd2901: y = 16'h5A5D;
            12'd2902: y = 16'h5A55;
            12'd2903: y = 16'h5A4D;
            12'd2904: y = 16'h5A45;
            12'd2905: y = 16'h5A3D;
            12'd2906: y = 16'h5A35;
            12'd2907: y = 16'h5A2D;
            12'd2908: y = 16'h5A25;
            12'd2909: y = 16'h5A1D;
            12'd2910: y = 16'h5A15;
            12'd2911: y = 16'h5A0E;
            12'd2912: y = 16'h5A06;
            12'd2913: y = 16'h59FE;
            12'd2914: y = 16'h59F6;
            12'd2915: y = 16'h59EE;
            12'd2916: y = 16'h59E6;
            12'd2917: y = 16'h59DE;
            12'd2918: y = 16'h59D6;
            12'd2919: y = 16'h59CE;
            12'd2920: y = 16'h59C6;
            12'd2921: y = 16'h59BF;
            12'd2922: y = 16'h59B7;
            12'd2923: y = 16'h59AF;
            12'd2924: y = 16'h59A7;
            12'd2925: y = 16'h599F;
            12'd2926: y = 16'h5997;
            12'd2927: y = 16'h5990;
            12'd2928: y = 16'h5988;
            12'd2929: y = 16'h5980;
            12'd2930: y = 16'h5978;
            12'd2931: y = 16'h5970;
            12'd2932: y = 16'h5968;
            12'd2933: y = 16'h5961;
            12'd2934: y = 16'h5959;
            12'd2935: y = 16'h5951;
            12'd2936: y = 16'h5949;
            12'd2937: y = 16'h5941;
            12'd2938: y = 16'h593A;
            12'd2939: y = 16'h5932;
            12'd2940: y = 16'h592A;
            12'd2941: y = 16'h5922;
            12'd2942: y = 16'h591B;
            12'd2943: y = 16'h5913;
            12'd2944: y = 16'h590B;
            12'd2945: y = 16'h5903;
            12'd2946: y = 16'h58FC;
            12'd2947: y = 16'h58F4;
            12'd2948: y = 16'h58EC;
            12'd2949: y = 16'h58E4;
            12'd2950: y = 16'h58DD;
            12'd2951: y = 16'h58D5;
            12'd2952: y = 16'h58CD;
            12'd2953: y = 16'h58C6;
            12'd2954: y = 16'h58BE;
            12'd2955: y = 16'h58B6;
            12'd2956: y = 16'h58AF;
            12'd2957: y = 16'h58A7;
            12'd2958: y = 16'h589F;
            12'd2959: y = 16'h5898;
            12'd2960: y = 16'h5890;
            12'd2961: y = 16'h5888;
            12'd2962: y = 16'h5881;
            12'd2963: y = 16'h5879;
            12'd2964: y = 16'h5871;
            12'd2965: y = 16'h586A;
            12'd2966: y = 16'h5862;
            12'd2967: y = 16'h585A;
            12'd2968: y = 16'h5853;
            12'd2969: y = 16'h584B;
            12'd2970: y = 16'h5844;
            12'd2971: y = 16'h583C;
            12'd2972: y = 16'h5834;
            12'd2973: y = 16'h582D;
            12'd2974: y = 16'h5825;
            12'd2975: y = 16'h581E;
            12'd2976: y = 16'h5816;
            12'd2977: y = 16'h580E;
            12'd2978: y = 16'h5807;
            12'd2979: y = 16'h57FF;
            12'd2980: y = 16'h57F8;
            12'd2981: y = 16'h57F0;
            12'd2982: y = 16'h57E9;
            12'd2983: y = 16'h57E1;
            12'd2984: y = 16'h57DA;
            12'd2985: y = 16'h57D2;
            12'd2986: y = 16'h57CB;
            12'd2987: y = 16'h57C3;
            12'd2988: y = 16'h57BB;
            12'd2989: y = 16'h57B4;
            12'd2990: y = 16'h57AC;
            12'd2991: y = 16'h57A5;
            12'd2992: y = 16'h579D;
            12'd2993: y = 16'h5796;
            12'd2994: y = 16'h578E;
            12'd2995: y = 16'h5787;
            12'd2996: y = 16'h577F;
            12'd2997: y = 16'h5778;
            12'd2998: y = 16'h5771;
            12'd2999: y = 16'h5769;
            12'd3000: y = 16'h5762;
            12'd3001: y = 16'h575A;
            12'd3002: y = 16'h5753;
            12'd3003: y = 16'h574B;
            12'd3004: y = 16'h5744;
            12'd3005: y = 16'h573C;
            12'd3006: y = 16'h5735;
            12'd3007: y = 16'h572E;
            12'd3008: y = 16'h5726;
            12'd3009: y = 16'h571F;
            12'd3010: y = 16'h5717;
            12'd3011: y = 16'h5710;
            12'd3012: y = 16'h5708;
            12'd3013: y = 16'h5701;
            12'd3014: y = 16'h56FA;
            12'd3015: y = 16'h56F2;
            12'd3016: y = 16'h56EB;
            12'd3017: y = 16'h56E4;
            12'd3018: y = 16'h56DC;
            12'd3019: y = 16'h56D5;
            12'd3020: y = 16'h56CD;
            12'd3021: y = 16'h56C6;
            12'd3022: y = 16'h56BF;
            12'd3023: y = 16'h56B7;
            12'd3024: y = 16'h56B0;
            12'd3025: y = 16'h56A9;
            12'd3026: y = 16'h56A1;
            12'd3027: y = 16'h569A;
            12'd3028: y = 16'h5693;
            12'd3029: y = 16'h568B;
            12'd3030: y = 16'h5684;
            12'd3031: y = 16'h567D;
            12'd3032: y = 16'h5676;
            12'd3033: y = 16'h566E;
            12'd3034: y = 16'h5667;
            12'd3035: y = 16'h5660;
            12'd3036: y = 16'h5658;
            12'd3037: y = 16'h5651;
            12'd3038: y = 16'h564A;
            12'd3039: y = 16'h5643;
            12'd3040: y = 16'h563B;
            12'd3041: y = 16'h5634;
            12'd3042: y = 16'h562D;
            12'd3043: y = 16'h5626;
            12'd3044: y = 16'h561E;
            12'd3045: y = 16'h5617;
            12'd3046: y = 16'h5610;
            12'd3047: y = 16'h5609;
            12'd3048: y = 16'h5601;
            12'd3049: y = 16'h55FA;
            12'd3050: y = 16'h55F3;
            12'd3051: y = 16'h55EC;
            12'd3052: y = 16'h55E4;
            12'd3053: y = 16'h55DD;
            12'd3054: y = 16'h55D6;
            12'd3055: y = 16'h55CF;
            12'd3056: y = 16'h55C8;
            12'd3057: y = 16'h55C1;
            12'd3058: y = 16'h55B9;
            12'd3059: y = 16'h55B2;
            12'd3060: y = 16'h55AB;
            12'd3061: y = 16'h55A4;
            12'd3062: y = 16'h559D;
            12'd3063: y = 16'h5596;
            12'd3064: y = 16'h558E;
            12'd3065: y = 16'h5587;
            12'd3066: y = 16'h5580;
            12'd3067: y = 16'h5579;
            12'd3068: y = 16'h5572;
            12'd3069: y = 16'h556B;
            12'd3070: y = 16'h5564;
            12'd3071: y = 16'h555C;
            12'd3072: y = 16'h5555;
            12'd3073: y = 16'h554E;
            12'd3074: y = 16'h5547;
            12'd3075: y = 16'h5540;
            12'd3076: y = 16'h5539;
            12'd3077: y = 16'h5532;
            12'd3078: y = 16'h552B;
            12'd3079: y = 16'h5524;
            12'd3080: y = 16'h551D;
            12'd3081: y = 16'h5516;
            12'd3082: y = 16'h550E;
            12'd3083: y = 16'h5507;
            12'd3084: y = 16'h5500;
            12'd3085: y = 16'h54F9;
            12'd3086: y = 16'h54F2;
            12'd3087: y = 16'h54EB;
            12'd3088: y = 16'h54E4;
            12'd3089: y = 16'h54DD;
            12'd3090: y = 16'h54D6;
            12'd3091: y = 16'h54CF;
            12'd3092: y = 16'h54C8;
            12'd3093: y = 16'h54C1;
            12'd3094: y = 16'h54BA;
            12'd3095: y = 16'h54B3;
            12'd3096: y = 16'h54AC;
            12'd3097: y = 16'h54A5;
            12'd3098: y = 16'h549E;
            12'd3099: y = 16'h5497;
            12'd3100: y = 16'h5490;
            12'd3101: y = 16'h5489;
            12'd3102: y = 16'h5482;
            12'd3103: y = 16'h547B;
            12'd3104: y = 16'h5474;
            12'd3105: y = 16'h546D;
            12'd3106: y = 16'h5466;
            12'd3107: y = 16'h545F;
            12'd3108: y = 16'h5458;
            12'd3109: y = 16'h5451;
            12'd3110: y = 16'h544A;
            12'd3111: y = 16'h5443;
            12'd3112: y = 16'h543D;
            12'd3113: y = 16'h5436;
            12'd3114: y = 16'h542F;
            12'd3115: y = 16'h5428;
            12'd3116: y = 16'h5421;
            12'd3117: y = 16'h541A;
            12'd3118: y = 16'h5413;
            12'd3119: y = 16'h540C;
            12'd3120: y = 16'h5405;
            12'd3121: y = 16'h53FE;
            12'd3122: y = 16'h53F7;
            12'd3123: y = 16'h53F1;
            12'd3124: y = 16'h53EA;
            12'd3125: y = 16'h53E3;
            12'd3126: y = 16'h53DC;
            12'd3127: y = 16'h53D5;
            12'd3128: y = 16'h53CE;
            12'd3129: y = 16'h53C7;
            12'd3130: y = 16'h53C1;
            12'd3131: y = 16'h53BA;
            12'd3132: y = 16'h53B3;
            12'd3133: y = 16'h53AC;
            12'd3134: y = 16'h53A5;
            12'd3135: y = 16'h539E;
            12'd3136: y = 16'h5398;
            12'd3137: y = 16'h5391;
            12'd3138: y = 16'h538A;
            12'd3139: y = 16'h5383;
            12'd3140: y = 16'h537C;
            12'd3141: y = 16'h5375;
            12'd3142: y = 16'h536F;
            12'd3143: y = 16'h5368;
            12'd3144: y = 16'h5361;
            12'd3145: y = 16'h535A;
            12'd3146: y = 16'h5353;
            12'd3147: y = 16'h534D;
            12'd3148: y = 16'h5346;
            12'd3149: y = 16'h533F;
            12'd3150: y = 16'h5338;
            12'd3151: y = 16'h5332;
            12'd3152: y = 16'h532B;
            12'd3153: y = 16'h5324;
            12'd3154: y = 16'h531D;
            12'd3155: y = 16'h5317;
            12'd3156: y = 16'h5310;
            12'd3157: y = 16'h5309;
            12'd3158: y = 16'h5302;
            12'd3159: y = 16'h52FC;
            12'd3160: y = 16'h52F5;
            12'd3161: y = 16'h52EE;
            12'd3162: y = 16'h52E8;
            12'd3163: y = 16'h52E1;
            12'd3164: y = 16'h52DA;
            12'd3165: y = 16'h52D3;
            12'd3166: y = 16'h52CD;
            12'd3167: y = 16'h52C6;
            12'd3168: y = 16'h52BF;
            12'd3169: y = 16'h52B9;
            12'd3170: y = 16'h52B2;
            12'd3171: y = 16'h52AB;
            12'd3172: y = 16'h52A5;
            12'd3173: y = 16'h529E;
            12'd3174: y = 16'h5297;
            12'd3175: y = 16'h5291;
            12'd3176: y = 16'h528A;
            12'd3177: y = 16'h5283;
            12'd3178: y = 16'h527D;
            12'd3179: y = 16'h5276;
            12'd3180: y = 16'h526F;
            12'd3181: y = 16'h5269;
            12'd3182: y = 16'h5262;
            12'd3183: y = 16'h525C;
            12'd3184: y = 16'h5255;
            12'd3185: y = 16'h524E;
            12'd3186: y = 16'h5248;
            12'd3187: y = 16'h5241;
            12'd3188: y = 16'h523A;
            12'd3189: y = 16'h5234;
            12'd3190: y = 16'h522D;
            12'd3191: y = 16'h5227;
            12'd3192: y = 16'h5220;
            12'd3193: y = 16'h5219;
            12'd3194: y = 16'h5213;
            12'd3195: y = 16'h520C;
            12'd3196: y = 16'h5206;
            12'd3197: y = 16'h51FF;
            12'd3198: y = 16'h51F9;
            12'd3199: y = 16'h51F2;
            12'd3200: y = 16'h51EC;
            12'd3201: y = 16'h51E5;
            12'd3202: y = 16'h51DE;
            12'd3203: y = 16'h51D8;
            12'd3204: y = 16'h51D1;
            12'd3205: y = 16'h51CB;
            12'd3206: y = 16'h51C4;
            12'd3207: y = 16'h51BE;
            12'd3208: y = 16'h51B7;
            12'd3209: y = 16'h51B1;
            12'd3210: y = 16'h51AA;
            12'd3211: y = 16'h51A4;
            12'd3212: y = 16'h519D;
            12'd3213: y = 16'h5197;
            12'd3214: y = 16'h5190;
            12'd3215: y = 16'h518A;
            12'd3216: y = 16'h5183;
            12'd3217: y = 16'h517D;
            12'd3218: y = 16'h5176;
            12'd3219: y = 16'h5170;
            12'd3220: y = 16'h5169;
            12'd3221: y = 16'h5163;
            12'd3222: y = 16'h515C;
            12'd3223: y = 16'h5156;
            12'd3224: y = 16'h514F;
            12'd3225: y = 16'h5149;
            12'd3226: y = 16'h5142;
            12'd3227: y = 16'h513C;
            12'd3228: y = 16'h5136;
            12'd3229: y = 16'h512F;
            12'd3230: y = 16'h5129;
            12'd3231: y = 16'h5122;
            12'd3232: y = 16'h511C;
            12'd3233: y = 16'h5115;
            12'd3234: y = 16'h510F;
            12'd3235: y = 16'h5109;
            12'd3236: y = 16'h5102;
            12'd3237: y = 16'h50FC;
            12'd3238: y = 16'h50F5;
            12'd3239: y = 16'h50EF;
            12'd3240: y = 16'h50E9;
            12'd3241: y = 16'h50E2;
            12'd3242: y = 16'h50DC;
            12'd3243: y = 16'h50D5;
            12'd3244: y = 16'h50CF;
            12'd3245: y = 16'h50C9;
            12'd3246: y = 16'h50C2;
            12'd3247: y = 16'h50BC;
            12'd3248: y = 16'h50B6;
            12'd3249: y = 16'h50AF;
            12'd3250: y = 16'h50A9;
            12'd3251: y = 16'h50A3;
            12'd3252: y = 16'h509C;
            12'd3253: y = 16'h5096;
            12'd3254: y = 16'h508F;
            12'd3255: y = 16'h5089;
            12'd3256: y = 16'h5083;
            12'd3257: y = 16'h507D;
            12'd3258: y = 16'h5076;
            12'd3259: y = 16'h5070;
            12'd3260: y = 16'h506A;
            12'd3261: y = 16'h5063;
            12'd3262: y = 16'h505D;
            12'd3263: y = 16'h5057;
            12'd3264: y = 16'h5050;
            12'd3265: y = 16'h504A;
            12'd3266: y = 16'h5044;
            12'd3267: y = 16'h503D;
            12'd3268: y = 16'h5037;
            12'd3269: y = 16'h5031;
            12'd3270: y = 16'h502B;
            12'd3271: y = 16'h5024;
            12'd3272: y = 16'h501E;
            12'd3273: y = 16'h5018;
            12'd3274: y = 16'h5012;
            12'd3275: y = 16'h500B;
            12'd3276: y = 16'h5005;
            12'd3277: y = 16'h4FFF;
            12'd3278: y = 16'h4FF9;
            12'd3279: y = 16'h4FF2;
            12'd3280: y = 16'h4FEC;
            12'd3281: y = 16'h4FE6;
            12'd3282: y = 16'h4FE0;
            12'd3283: y = 16'h4FD9;
            12'd3284: y = 16'h4FD3;
            12'd3285: y = 16'h4FCD;
            12'd3286: y = 16'h4FC7;
            12'd3287: y = 16'h4FC0;
            12'd3288: y = 16'h4FBA;
            12'd3289: y = 16'h4FB4;
            12'd3290: y = 16'h4FAE;
            12'd3291: y = 16'h4FA8;
            12'd3292: y = 16'h4FA1;
            12'd3293: y = 16'h4F9B;
            12'd3294: y = 16'h4F95;
            12'd3295: y = 16'h4F8F;
            12'd3296: y = 16'h4F89;
            12'd3297: y = 16'h4F83;
            12'd3298: y = 16'h4F7C;
            12'd3299: y = 16'h4F76;
            12'd3300: y = 16'h4F70;
            12'd3301: y = 16'h4F6A;
            12'd3302: y = 16'h4F64;
            12'd3303: y = 16'h4F5E;
            12'd3304: y = 16'h4F57;
            12'd3305: y = 16'h4F51;
            12'd3306: y = 16'h4F4B;
            12'd3307: y = 16'h4F45;
            12'd3308: y = 16'h4F3F;
            12'd3309: y = 16'h4F39;
            12'd3310: y = 16'h4F33;
            12'd3311: y = 16'h4F2C;
            12'd3312: y = 16'h4F26;
            12'd3313: y = 16'h4F20;
            12'd3314: y = 16'h4F1A;
            12'd3315: y = 16'h4F14;
            12'd3316: y = 16'h4F0E;
            12'd3317: y = 16'h4F08;
            12'd3318: y = 16'h4F02;
            12'd3319: y = 16'h4EFC;
            12'd3320: y = 16'h4EF6;
            12'd3321: y = 16'h4EEF;
            12'd3322: y = 16'h4EE9;
            12'd3323: y = 16'h4EE3;
            12'd3324: y = 16'h4EDD;
            12'd3325: y = 16'h4ED7;
            12'd3326: y = 16'h4ED1;
            12'd3327: y = 16'h4ECB;
            12'd3328: y = 16'h4EC5;
            12'd3329: y = 16'h4EBF;
            12'd3330: y = 16'h4EB9;
            12'd3331: y = 16'h4EB3;
            12'd3332: y = 16'h4EAD;
            12'd3333: y = 16'h4EA7;
            12'd3334: y = 16'h4EA1;
            12'd3335: y = 16'h4E9B;
            12'd3336: y = 16'h4E95;
            12'd3337: y = 16'h4E8F;
            12'd3338: y = 16'h4E89;
            12'd3339: y = 16'h4E82;
            12'd3340: y = 16'h4E7C;
            12'd3341: y = 16'h4E76;
            12'd3342: y = 16'h4E70;
            12'd3343: y = 16'h4E6A;
            12'd3344: y = 16'h4E64;
            12'd3345: y = 16'h4E5E;
            12'd3346: y = 16'h4E58;
            12'd3347: y = 16'h4E52;
            12'd3348: y = 16'h4E4C;
            12'd3349: y = 16'h4E46;
            12'd3350: y = 16'h4E40;
            12'd3351: y = 16'h4E3B;
            12'd3352: y = 16'h4E35;
            12'd3353: y = 16'h4E2F;
            12'd3354: y = 16'h4E29;
            12'd3355: y = 16'h4E23;
            12'd3356: y = 16'h4E1D;
            12'd3357: y = 16'h4E17;
            12'd3358: y = 16'h4E11;
            12'd3359: y = 16'h4E0B;
            12'd3360: y = 16'h4E05;
            12'd3361: y = 16'h4DFF;
            12'd3362: y = 16'h4DF9;
            12'd3363: y = 16'h4DF3;
            12'd3364: y = 16'h4DED;
            12'd3365: y = 16'h4DE7;
            12'd3366: y = 16'h4DE1;
            12'd3367: y = 16'h4DDB;
            12'd3368: y = 16'h4DD5;
            12'd3369: y = 16'h4DD0;
            12'd3370: y = 16'h4DCA;
            12'd3371: y = 16'h4DC4;
            12'd3372: y = 16'h4DBE;
            12'd3373: y = 16'h4DB8;
            12'd3374: y = 16'h4DB2;
            12'd3375: y = 16'h4DAC;
            12'd3376: y = 16'h4DA6;
            12'd3377: y = 16'h4DA0;
            12'd3378: y = 16'h4D9A;
            12'd3379: y = 16'h4D95;
            12'd3380: y = 16'h4D8F;
            12'd3381: y = 16'h4D89;
            12'd3382: y = 16'h4D83;
            12'd3383: y = 16'h4D7D;
            12'd3384: y = 16'h4D77;
            12'd3385: y = 16'h4D71;
            12'd3386: y = 16'h4D6C;
            12'd3387: y = 16'h4D66;
            12'd3388: y = 16'h4D60;
            12'd3389: y = 16'h4D5A;
            12'd3390: y = 16'h4D54;
            12'd3391: y = 16'h4D4E;
            12'd3392: y = 16'h4D48;
            12'd3393: y = 16'h4D43;
            12'd3394: y = 16'h4D3D;
            12'd3395: y = 16'h4D37;
            12'd3396: y = 16'h4D31;
            12'd3397: y = 16'h4D2B;
            12'd3398: y = 16'h4D26;
            12'd3399: y = 16'h4D20;
            12'd3400: y = 16'h4D1A;
            12'd3401: y = 16'h4D14;
            12'd3402: y = 16'h4D0E;
            12'd3403: y = 16'h4D09;
            12'd3404: y = 16'h4D03;
            12'd3405: y = 16'h4CFD;
            12'd3406: y = 16'h4CF7;
            12'd3407: y = 16'h4CF1;
            12'd3408: y = 16'h4CEC;
            12'd3409: y = 16'h4CE6;
            12'd3410: y = 16'h4CE0;
            12'd3411: y = 16'h4CDA;
            12'd3412: y = 16'h4CD4;
            12'd3413: y = 16'h4CCF;
            12'd3414: y = 16'h4CC9;
            12'd3415: y = 16'h4CC3;
            12'd3416: y = 16'h4CBD;
            12'd3417: y = 16'h4CB8;
            12'd3418: y = 16'h4CB2;
            12'd3419: y = 16'h4CAC;
            12'd3420: y = 16'h4CA6;
            12'd3421: y = 16'h4CA1;
            12'd3422: y = 16'h4C9B;
            12'd3423: y = 16'h4C95;
            12'd3424: y = 16'h4C90;
            12'd3425: y = 16'h4C8A;
            12'd3426: y = 16'h4C84;
            12'd3427: y = 16'h4C7E;
            12'd3428: y = 16'h4C79;
            12'd3429: y = 16'h4C73;
            12'd3430: y = 16'h4C6D;
            12'd3431: y = 16'h4C68;
            12'd3432: y = 16'h4C62;
            12'd3433: y = 16'h4C5C;
            12'd3434: y = 16'h4C56;
            12'd3435: y = 16'h4C51;
            12'd3436: y = 16'h4C4B;
            12'd3437: y = 16'h4C45;
            12'd3438: y = 16'h4C40;
            12'd3439: y = 16'h4C3A;
            12'd3440: y = 16'h4C34;
            12'd3441: y = 16'h4C2F;
            12'd3442: y = 16'h4C29;
            12'd3443: y = 16'h4C23;
            12'd3444: y = 16'h4C1E;
            12'd3445: y = 16'h4C18;
            12'd3446: y = 16'h4C12;
            12'd3447: y = 16'h4C0D;
            12'd3448: y = 16'h4C07;
            12'd3449: y = 16'h4C01;
            12'd3450: y = 16'h4BFC;
            12'd3451: y = 16'h4BF6;
            12'd3452: y = 16'h4BF1;
            12'd3453: y = 16'h4BEB;
            12'd3454: y = 16'h4BE5;
            12'd3455: y = 16'h4BE0;
            12'd3456: y = 16'h4BDA;
            12'd3457: y = 16'h4BD4;
            12'd3458: y = 16'h4BCF;
            12'd3459: y = 16'h4BC9;
            12'd3460: y = 16'h4BC4;
            12'd3461: y = 16'h4BBE;
            12'd3462: y = 16'h4BB8;
            12'd3463: y = 16'h4BB3;
            12'd3464: y = 16'h4BAD;
            12'd3465: y = 16'h4BA8;
            12'd3466: y = 16'h4BA2;
            12'd3467: y = 16'h4B9C;
            12'd3468: y = 16'h4B97;
            12'd3469: y = 16'h4B91;
            12'd3470: y = 16'h4B8C;
            12'd3471: y = 16'h4B86;
            12'd3472: y = 16'h4B81;
            12'd3473: y = 16'h4B7B;
            12'd3474: y = 16'h4B75;
            12'd3475: y = 16'h4B70;
            12'd3476: y = 16'h4B6A;
            12'd3477: y = 16'h4B65;
            12'd3478: y = 16'h4B5F;
            12'd3479: y = 16'h4B5A;
            12'd3480: y = 16'h4B54;
            12'd3481: y = 16'h4B4F;
            12'd3482: y = 16'h4B49;
            12'd3483: y = 16'h4B44;
            12'd3484: y = 16'h4B3E;
            12'd3485: y = 16'h4B38;
            12'd3486: y = 16'h4B33;
            12'd3487: y = 16'h4B2D;
            12'd3488: y = 16'h4B28;
            12'd3489: y = 16'h4B22;
            12'd3490: y = 16'h4B1D;
            12'd3491: y = 16'h4B17;
            12'd3492: y = 16'h4B12;
            12'd3493: y = 16'h4B0C;
            12'd3494: y = 16'h4B07;
            12'd3495: y = 16'h4B01;
            12'd3496: y = 16'h4AFC;
            12'd3497: y = 16'h4AF6;
            12'd3498: y = 16'h4AF1;
            12'd3499: y = 16'h4AEB;
            12'd3500: y = 16'h4AE6;
            12'd3501: y = 16'h4AE0;
            12'd3502: y = 16'h4ADB;
            12'd3503: y = 16'h4AD6;
            12'd3504: y = 16'h4AD0;
            12'd3505: y = 16'h4ACB;
            12'd3506: y = 16'h4AC5;
            12'd3507: y = 16'h4AC0;
            12'd3508: y = 16'h4ABA;
            12'd3509: y = 16'h4AB5;
            12'd3510: y = 16'h4AAF;
            12'd3511: y = 16'h4AAA;
            12'd3512: y = 16'h4AA4;
            12'd3513: y = 16'h4A9F;
            12'd3514: y = 16'h4A9A;
            12'd3515: y = 16'h4A94;
            12'd3516: y = 16'h4A8F;
            12'd3517: y = 16'h4A89;
            12'd3518: y = 16'h4A84;
            12'd3519: y = 16'h4A7E;
            12'd3520: y = 16'h4A79;
            12'd3521: y = 16'h4A74;
            12'd3522: y = 16'h4A6E;
            12'd3523: y = 16'h4A69;
            12'd3524: y = 16'h4A63;
            12'd3525: y = 16'h4A5E;
            12'd3526: y = 16'h4A59;
            12'd3527: y = 16'h4A53;
            12'd3528: y = 16'h4A4E;
            12'd3529: y = 16'h4A48;
            12'd3530: y = 16'h4A43;
            12'd3531: y = 16'h4A3E;
            12'd3532: y = 16'h4A38;
            12'd3533: y = 16'h4A33;
            12'd3534: y = 16'h4A2D;
            12'd3535: y = 16'h4A28;
            12'd3536: y = 16'h4A23;
            12'd3537: y = 16'h4A1D;
            12'd3538: y = 16'h4A18;
            12'd3539: y = 16'h4A13;
            12'd3540: y = 16'h4A0D;
            12'd3541: y = 16'h4A08;
            12'd3542: y = 16'h4A03;
            12'd3543: y = 16'h49FD;
            12'd3544: y = 16'h49F8;
            12'd3545: y = 16'h49F3;
            12'd3546: y = 16'h49ED;
            12'd3547: y = 16'h49E8;
            12'd3548: y = 16'h49E3;
            12'd3549: y = 16'h49DD;
            12'd3550: y = 16'h49D8;
            12'd3551: y = 16'h49D3;
            12'd3552: y = 16'h49CD;
            12'd3553: y = 16'h49C8;
            12'd3554: y = 16'h49C3;
            12'd3555: y = 16'h49BD;
            12'd3556: y = 16'h49B8;
            12'd3557: y = 16'h49B3;
            12'd3558: y = 16'h49AD;
            12'd3559: y = 16'h49A8;
            12'd3560: y = 16'h49A3;
            12'd3561: y = 16'h499E;
            12'd3562: y = 16'h4998;
            12'd3563: y = 16'h4993;
            12'd3564: y = 16'h498E;
            12'd3565: y = 16'h4988;
            12'd3566: y = 16'h4983;
            12'd3567: y = 16'h497E;
            12'd3568: y = 16'h4979;
            12'd3569: y = 16'h4973;
            12'd3570: y = 16'h496E;
            12'd3571: y = 16'h4969;
            12'd3572: y = 16'h4963;
            12'd3573: y = 16'h495E;
            12'd3574: y = 16'h4959;
            12'd3575: y = 16'h4954;
            12'd3576: y = 16'h494E;
            12'd3577: y = 16'h4949;
            12'd3578: y = 16'h4944;
            12'd3579: y = 16'h493F;
            12'd3580: y = 16'h4939;
            12'd3581: y = 16'h4934;
            12'd3582: y = 16'h492F;
            12'd3583: y = 16'h492A;
            12'd3584: y = 16'h4925;
            12'd3585: y = 16'h491F;
            12'd3586: y = 16'h491A;
            12'd3587: y = 16'h4915;
            12'd3588: y = 16'h4910;
            12'd3589: y = 16'h490A;
            12'd3590: y = 16'h4905;
            12'd3591: y = 16'h4900;
            12'd3592: y = 16'h48FB;
            12'd3593: y = 16'h48F6;
            12'd3594: y = 16'h48F0;
            12'd3595: y = 16'h48EB;
            12'd3596: y = 16'h48E6;
            12'd3597: y = 16'h48E1;
            12'd3598: y = 16'h48DC;
            12'd3599: y = 16'h48D7;
            12'd3600: y = 16'h48D1;
            12'd3601: y = 16'h48CC;
            12'd3602: y = 16'h48C7;
            12'd3603: y = 16'h48C2;
            12'd3604: y = 16'h48BD;
            12'd3605: y = 16'h48B7;
            12'd3606: y = 16'h48B2;
            12'd3607: y = 16'h48AD;
            12'd3608: y = 16'h48A8;
            12'd3609: y = 16'h48A3;
            12'd3610: y = 16'h489E;
            12'd3611: y = 16'h4899;
            12'd3612: y = 16'h4893;
            12'd3613: y = 16'h488E;
            12'd3614: y = 16'h4889;
            12'd3615: y = 16'h4884;
            12'd3616: y = 16'h487F;
            12'd3617: y = 16'h487A;
            12'd3618: y = 16'h4875;
            12'd3619: y = 16'h486F;
            12'd3620: y = 16'h486A;
            12'd3621: y = 16'h4865;
            12'd3622: y = 16'h4860;
            12'd3623: y = 16'h485B;
            12'd3624: y = 16'h4856;
            12'd3625: y = 16'h4851;
            12'd3626: y = 16'h484C;
            12'd3627: y = 16'h4847;
            12'd3628: y = 16'h4841;
            12'd3629: y = 16'h483C;
            12'd3630: y = 16'h4837;
            12'd3631: y = 16'h4832;
            12'd3632: y = 16'h482D;
            12'd3633: y = 16'h4828;
            12'd3634: y = 16'h4823;
            12'd3635: y = 16'h481E;
            12'd3636: y = 16'h4819;
            12'd3637: y = 16'h4814;
            12'd3638: y = 16'h480F;
            12'd3639: y = 16'h480A;
            12'd3640: y = 16'h4805;
            12'd3641: y = 16'h47FF;
            12'd3642: y = 16'h47FA;
            12'd3643: y = 16'h47F5;
            12'd3644: y = 16'h47F0;
            12'd3645: y = 16'h47EB;
            12'd3646: y = 16'h47E6;
            12'd3647: y = 16'h47E1;
            12'd3648: y = 16'h47DC;
            12'd3649: y = 16'h47D7;
            12'd3650: y = 16'h47D2;
            12'd3651: y = 16'h47CD;
            12'd3652: y = 16'h47C8;
            12'd3653: y = 16'h47C3;
            12'd3654: y = 16'h47BE;
            12'd3655: y = 16'h47B9;
            12'd3656: y = 16'h47B4;
            12'd3657: y = 16'h47AF;
            12'd3658: y = 16'h47AA;
            12'd3659: y = 16'h47A5;
            12'd3660: y = 16'h47A0;
            12'd3661: y = 16'h479B;
            12'd3662: y = 16'h4796;
            12'd3663: y = 16'h4791;
            12'd3664: y = 16'h478C;
            12'd3665: y = 16'h4787;
            12'd3666: y = 16'h4782;
            12'd3667: y = 16'h477D;
            12'd3668: y = 16'h4778;
            12'd3669: y = 16'h4773;
            12'd3670: y = 16'h476E;
            12'd3671: y = 16'h4769;
            12'd3672: y = 16'h4764;
            12'd3673: y = 16'h475F;
            12'd3674: y = 16'h475A;
            12'd3675: y = 16'h4755;
            12'd3676: y = 16'h4750;
            12'd3677: y = 16'h474B;
            12'd3678: y = 16'h4746;
            12'd3679: y = 16'h4741;
            12'd3680: y = 16'h473C;
            12'd3681: y = 16'h4737;
            12'd3682: y = 16'h4732;
            12'd3683: y = 16'h472D;
            12'd3684: y = 16'h4728;
            12'd3685: y = 16'h4723;
            12'd3686: y = 16'h471E;
            12'd3687: y = 16'h4719;
            12'd3688: y = 16'h4715;
            12'd3689: y = 16'h4710;
            12'd3690: y = 16'h470B;
            12'd3691: y = 16'h4706;
            12'd3692: y = 16'h4701;
            12'd3693: y = 16'h46FC;
            12'd3694: y = 16'h46F7;
            12'd3695: y = 16'h46F2;
            12'd3696: y = 16'h46ED;
            12'd3697: y = 16'h46E8;
            12'd3698: y = 16'h46E3;
            12'd3699: y = 16'h46DE;
            12'd3700: y = 16'h46DA;
            12'd3701: y = 16'h46D5;
            12'd3702: y = 16'h46D0;
            12'd3703: y = 16'h46CB;
            12'd3704: y = 16'h46C6;
            12'd3705: y = 16'h46C1;
            12'd3706: y = 16'h46BC;
            12'd3707: y = 16'h46B7;
            12'd3708: y = 16'h46B2;
            12'd3709: y = 16'h46AE;
            12'd3710: y = 16'h46A9;
            12'd3711: y = 16'h46A4;
            12'd3712: y = 16'h469F;
            12'd3713: y = 16'h469A;
            12'd3714: y = 16'h4695;
            12'd3715: y = 16'h4690;
            12'd3716: y = 16'h468B;
            12'd3717: y = 16'h4687;
            12'd3718: y = 16'h4682;
            12'd3719: y = 16'h467D;
            12'd3720: y = 16'h4678;
            12'd3721: y = 16'h4673;
            12'd3722: y = 16'h466E;
            12'd3723: y = 16'h4669;
            12'd3724: y = 16'h4665;
            12'd3725: y = 16'h4660;
            12'd3726: y = 16'h465B;
            12'd3727: y = 16'h4656;
            12'd3728: y = 16'h4651;
            12'd3729: y = 16'h464C;
            12'd3730: y = 16'h4648;
            12'd3731: y = 16'h4643;
            12'd3732: y = 16'h463E;
            12'd3733: y = 16'h4639;
            12'd3734: y = 16'h4634;
            12'd3735: y = 16'h4630;
            12'd3736: y = 16'h462B;
            12'd3737: y = 16'h4626;
            12'd3738: y = 16'h4621;
            12'd3739: y = 16'h461C;
            12'd3740: y = 16'h4618;
            12'd3741: y = 16'h4613;
            12'd3742: y = 16'h460E;
            12'd3743: y = 16'h4609;
            12'd3744: y = 16'h4604;
            12'd3745: y = 16'h4600;
            12'd3746: y = 16'h45FB;
            12'd3747: y = 16'h45F6;
            12'd3748: y = 16'h45F1;
            12'd3749: y = 16'h45EC;
            12'd3750: y = 16'h45E8;
            12'd3751: y = 16'h45E3;
            12'd3752: y = 16'h45DE;
            12'd3753: y = 16'h45D9;
            12'd3754: y = 16'h45D5;
            12'd3755: y = 16'h45D0;
            12'd3756: y = 16'h45CB;
            12'd3757: y = 16'h45C6;
            12'd3758: y = 16'h45C2;
            12'd3759: y = 16'h45BD;
            12'd3760: y = 16'h45B8;
            12'd3761: y = 16'h45B3;
            12'd3762: y = 16'h45AF;
            12'd3763: y = 16'h45AA;
            12'd3764: y = 16'h45A5;
            12'd3765: y = 16'h45A0;
            12'd3766: y = 16'h459C;
            12'd3767: y = 16'h4597;
            12'd3768: y = 16'h4592;
            12'd3769: y = 16'h458D;
            12'd3770: y = 16'h4589;
            12'd3771: y = 16'h4584;
            12'd3772: y = 16'h457F;
            12'd3773: y = 16'h457B;
            12'd3774: y = 16'h4576;
            12'd3775: y = 16'h4571;
            12'd3776: y = 16'h456C;
            12'd3777: y = 16'h4568;
            12'd3778: y = 16'h4563;
            12'd3779: y = 16'h455E;
            12'd3780: y = 16'h455A;
            12'd3781: y = 16'h4555;
            12'd3782: y = 16'h4550;
            12'd3783: y = 16'h454C;
            12'd3784: y = 16'h4547;
            12'd3785: y = 16'h4542;
            12'd3786: y = 16'h453E;
            12'd3787: y = 16'h4539;
            12'd3788: y = 16'h4534;
            12'd3789: y = 16'h452F;
            12'd3790: y = 16'h452B;
            12'd3791: y = 16'h4526;
            12'd3792: y = 16'h4521;
            12'd3793: y = 16'h451D;
            12'd3794: y = 16'h4518;
            12'd3795: y = 16'h4513;
            12'd3796: y = 16'h450F;
            12'd3797: y = 16'h450A;
            12'd3798: y = 16'h4506;
            12'd3799: y = 16'h4501;
            12'd3800: y = 16'h44FC;
            12'd3801: y = 16'h44F8;
            12'd3802: y = 16'h44F3;
            12'd3803: y = 16'h44EE;
            12'd3804: y = 16'h44EA;
            12'd3805: y = 16'h44E5;
            12'd3806: y = 16'h44E0;
            12'd3807: y = 16'h44DC;
            12'd3808: y = 16'h44D7;
            12'd3809: y = 16'h44D2;
            12'd3810: y = 16'h44CE;
            12'd3811: y = 16'h44C9;
            12'd3812: y = 16'h44C5;
            12'd3813: y = 16'h44C0;
            12'd3814: y = 16'h44BB;
            12'd3815: y = 16'h44B7;
            12'd3816: y = 16'h44B2;
            12'd3817: y = 16'h44AE;
            12'd3818: y = 16'h44A9;
            12'd3819: y = 16'h44A4;
            12'd3820: y = 16'h44A0;
            12'd3821: y = 16'h449B;
            12'd3822: y = 16'h4497;
            12'd3823: y = 16'h4492;
            12'd3824: y = 16'h448D;
            12'd3825: y = 16'h4489;
            12'd3826: y = 16'h4484;
            12'd3827: y = 16'h4480;
            12'd3828: y = 16'h447B;
            12'd3829: y = 16'h4476;
            12'd3830: y = 16'h4472;
            12'd3831: y = 16'h446D;
            12'd3832: y = 16'h4469;
            12'd3833: y = 16'h4464;
            12'd3834: y = 16'h4460;
            12'd3835: y = 16'h445B;
            12'd3836: y = 16'h4456;
            12'd3837: y = 16'h4452;
            12'd3838: y = 16'h444D;
            12'd3839: y = 16'h4449;
            12'd3840: y = 16'h4444;
            12'd3841: y = 16'h4440;
            12'd3842: y = 16'h443B;
            12'd3843: y = 16'h4437;
            12'd3844: y = 16'h4432;
            12'd3845: y = 16'h442E;
            12'd3846: y = 16'h4429;
            12'd3847: y = 16'h4424;
            12'd3848: y = 16'h4420;
            12'd3849: y = 16'h441B;
            12'd3850: y = 16'h4417;
            12'd3851: y = 16'h4412;
            12'd3852: y = 16'h440E;
            12'd3853: y = 16'h4409;
            12'd3854: y = 16'h4405;
            12'd3855: y = 16'h4400;
            12'd3856: y = 16'h43FC;
            12'd3857: y = 16'h43F7;
            12'd3858: y = 16'h43F3;
            12'd3859: y = 16'h43EE;
            12'd3860: y = 16'h43EA;
            12'd3861: y = 16'h43E5;
            12'd3862: y = 16'h43E1;
            12'd3863: y = 16'h43DC;
            12'd3864: y = 16'h43D8;
            12'd3865: y = 16'h43D3;
            12'd3866: y = 16'h43CF;
            12'd3867: y = 16'h43CA;
            12'd3868: y = 16'h43C6;
            12'd3869: y = 16'h43C1;
            12'd3870: y = 16'h43BD;
            12'd3871: y = 16'h43B8;
            12'd3872: y = 16'h43B4;
            12'd3873: y = 16'h43AF;
            12'd3874: y = 16'h43AB;
            12'd3875: y = 16'h43A6;
            12'd3876: y = 16'h43A2;
            12'd3877: y = 16'h439D;
            12'd3878: y = 16'h4399;
            12'd3879: y = 16'h4395;
            12'd3880: y = 16'h4390;
            12'd3881: y = 16'h438C;
            12'd3882: y = 16'h4387;
            12'd3883: y = 16'h4383;
            12'd3884: y = 16'h437E;
            12'd3885: y = 16'h437A;
            12'd3886: y = 16'h4375;
            12'd3887: y = 16'h4371;
            12'd3888: y = 16'h436D;
            12'd3889: y = 16'h4368;
            12'd3890: y = 16'h4364;
            12'd3891: y = 16'h435F;
            12'd3892: y = 16'h435B;
            12'd3893: y = 16'h4356;
            12'd3894: y = 16'h4352;
            12'd3895: y = 16'h434D;
            12'd3896: y = 16'h4349;
            12'd3897: y = 16'h4345;
            12'd3898: y = 16'h4340;
            12'd3899: y = 16'h433C;
            12'd3900: y = 16'h4337;
            12'd3901: y = 16'h4333;
            12'd3902: y = 16'h432F;
            12'd3903: y = 16'h432A;
            12'd3904: y = 16'h4326;
            12'd3905: y = 16'h4321;
            12'd3906: y = 16'h431D;
            12'd3907: y = 16'h4319;
            12'd3908: y = 16'h4314;
            12'd3909: y = 16'h4310;
            12'd3910: y = 16'h430B;
            12'd3911: y = 16'h4307;
            12'd3912: y = 16'h4303;
            12'd3913: y = 16'h42FE;
            12'd3914: y = 16'h42FA;
            12'd3915: y = 16'h42F5;
            12'd3916: y = 16'h42F1;
            12'd3917: y = 16'h42ED;
            12'd3918: y = 16'h42E8;
            12'd3919: y = 16'h42E4;
            12'd3920: y = 16'h42E0;
            12'd3921: y = 16'h42DB;
            12'd3922: y = 16'h42D7;
            12'd3923: y = 16'h42D3;
            12'd3924: y = 16'h42CE;
            12'd3925: y = 16'h42CA;
            12'd3926: y = 16'h42C5;
            12'd3927: y = 16'h42C1;
            12'd3928: y = 16'h42BD;
            12'd3929: y = 16'h42B8;
            12'd3930: y = 16'h42B4;
            12'd3931: y = 16'h42B0;
            12'd3932: y = 16'h42AB;
            12'd3933: y = 16'h42A7;
            12'd3934: y = 16'h42A3;
            12'd3935: y = 16'h429E;
            12'd3936: y = 16'h429A;
            12'd3937: y = 16'h4296;
            12'd3938: y = 16'h4291;
            12'd3939: y = 16'h428D;
            12'd3940: y = 16'h4289;
            12'd3941: y = 16'h4284;
            12'd3942: y = 16'h4280;
            12'd3943: y = 16'h427C;
            12'd3944: y = 16'h4277;
            12'd3945: y = 16'h4273;
            12'd3946: y = 16'h426F;
            12'd3947: y = 16'h426A;
            12'd3948: y = 16'h4266;
            12'd3949: y = 16'h4262;
            12'd3950: y = 16'h425E;
            12'd3951: y = 16'h4259;
            12'd3952: y = 16'h4255;
            12'd3953: y = 16'h4251;
            12'd3954: y = 16'h424C;
            12'd3955: y = 16'h4248;
            12'd3956: y = 16'h4244;
            12'd3957: y = 16'h4240;
            12'd3958: y = 16'h423B;
            12'd3959: y = 16'h4237;
            12'd3960: y = 16'h4233;
            12'd3961: y = 16'h422E;
            12'd3962: y = 16'h422A;
            12'd3963: y = 16'h4226;
            12'd3964: y = 16'h4222;
            12'd3965: y = 16'h421D;
            12'd3966: y = 16'h4219;
            12'd3967: y = 16'h4215;
            12'd3968: y = 16'h4211;
            12'd3969: y = 16'h420C;
            12'd3970: y = 16'h4208;
            12'd3971: y = 16'h4204;
            12'd3972: y = 16'h41FF;
            12'd3973: y = 16'h41FB;
            12'd3974: y = 16'h41F7;
            12'd3975: y = 16'h41F3;
            12'd3976: y = 16'h41EE;
            12'd3977: y = 16'h41EA;
            12'd3978: y = 16'h41E6;
            12'd3979: y = 16'h41E2;
            12'd3980: y = 16'h41DE;
            12'd3981: y = 16'h41D9;
            12'd3982: y = 16'h41D5;
            12'd3983: y = 16'h41D1;
            12'd3984: y = 16'h41CD;
            12'd3985: y = 16'h41C8;
            12'd3986: y = 16'h41C4;
            12'd3987: y = 16'h41C0;
            12'd3988: y = 16'h41BC;
            12'd3989: y = 16'h41B7;
            12'd3990: y = 16'h41B3;
            12'd3991: y = 16'h41AF;
            12'd3992: y = 16'h41AB;
            12'd3993: y = 16'h41A7;
            12'd3994: y = 16'h41A2;
            12'd3995: y = 16'h419E;
            12'd3996: y = 16'h419A;
            12'd3997: y = 16'h4196;
            12'd3998: y = 16'h4192;
            12'd3999: y = 16'h418D;
            12'd4000: y = 16'h4189;
            12'd4001: y = 16'h4185;
            12'd4002: y = 16'h4181;
            12'd4003: y = 16'h417D;
            12'd4004: y = 16'h4178;
            12'd4005: y = 16'h4174;
            12'd4006: y = 16'h4170;
            12'd4007: y = 16'h416C;
            12'd4008: y = 16'h4168;
            12'd4009: y = 16'h4164;
            12'd4010: y = 16'h415F;
            12'd4011: y = 16'h415B;
            12'd4012: y = 16'h4157;
            12'd4013: y = 16'h4153;
            12'd4014: y = 16'h414F;
            12'd4015: y = 16'h414B;
            12'd4016: y = 16'h4146;
            12'd4017: y = 16'h4142;
            12'd4018: y = 16'h413E;
            12'd4019: y = 16'h413A;
            12'd4020: y = 16'h4136;
            12'd4021: y = 16'h4132;
            12'd4022: y = 16'h412D;
            12'd4023: y = 16'h4129;
            12'd4024: y = 16'h4125;
            12'd4025: y = 16'h4121;
            12'd4026: y = 16'h411D;
            12'd4027: y = 16'h4119;
            12'd4028: y = 16'h4115;
            12'd4029: y = 16'h4110;
            12'd4030: y = 16'h410C;
            12'd4031: y = 16'h4108;
            12'd4032: y = 16'h4104;
            12'd4033: y = 16'h4100;
            12'd4034: y = 16'h40FC;
            12'd4035: y = 16'h40F8;
            12'd4036: y = 16'h40F4;
            12'd4037: y = 16'h40EF;
            12'd4038: y = 16'h40EB;
            12'd4039: y = 16'h40E7;
            12'd4040: y = 16'h40E3;
            12'd4041: y = 16'h40DF;
            12'd4042: y = 16'h40DB;
            12'd4043: y = 16'h40D7;
            12'd4044: y = 16'h40D3;
            12'd4045: y = 16'h40CF;
            12'd4046: y = 16'h40CA;
            12'd4047: y = 16'h40C6;
            12'd4048: y = 16'h40C2;
            12'd4049: y = 16'h40BE;
            12'd4050: y = 16'h40BA;
            12'd4051: y = 16'h40B6;
            12'd4052: y = 16'h40B2;
            12'd4053: y = 16'h40AE;
            12'd4054: y = 16'h40AA;
            12'd4055: y = 16'h40A6;
            12'd4056: y = 16'h40A2;
            12'd4057: y = 16'h409D;
            12'd4058: y = 16'h4099;
            12'd4059: y = 16'h4095;
            12'd4060: y = 16'h4091;
            12'd4061: y = 16'h408D;
            12'd4062: y = 16'h4089;
            12'd4063: y = 16'h4085;
            12'd4064: y = 16'h4081;
            12'd4065: y = 16'h407D;
            12'd4066: y = 16'h4079;
            12'd4067: y = 16'h4075;
            12'd4068: y = 16'h4071;
            12'd4069: y = 16'h406D;
            12'd4070: y = 16'h4069;
            12'd4071: y = 16'h4065;
            12'd4072: y = 16'h4061;
            12'd4073: y = 16'h405D;
            12'd4074: y = 16'h4058;
            12'd4075: y = 16'h4054;
            12'd4076: y = 16'h4050;
            12'd4077: y = 16'h404C;
            12'd4078: y = 16'h4048;
            12'd4079: y = 16'h4044;
            12'd4080: y = 16'h4040;
            12'd4081: y = 16'h403C;
            12'd4082: y = 16'h4038;
            12'd4083: y = 16'h4034;
            12'd4084: y = 16'h4030;
            12'd4085: y = 16'h402C;
            12'd4086: y = 16'h4028;
            12'd4087: y = 16'h4024;
            12'd4088: y = 16'h4020;
            12'd4089: y = 16'h401C;
            12'd4090: y = 16'h4018;
            12'd4091: y = 16'h4014;
            12'd4092: y = 16'h4010;
            12'd4093: y = 16'h400C;
            12'd4094: y = 16'h4008;
            12'd4095: y = 16'h4004;
            default:  y = 16'h0000;
        endcase
    end
endmodule
