module Transmission_Reciprocal_LUT (
    input      [15:0] in,  // Q0.16 Transmission value input (unsigned)
    output reg [15:0] out  // Q2.14 Inverse Transmission value output (unsigned)
);

    wire [11:0] scaled_in = in[15:4];
    
    always @(*) begin
        casez(scaled_in)
            12'd   0: out = 16'h4000;
            12'd   1: out = 16'hFFFF;
            12'd   2: out = 16'hFFFF;
            12'd   3: out = 16'hFFFF;
            12'd   4: out = 16'hFFFF;
            12'd   5: out = 16'hFFFF;
            12'd   6: out = 16'hFFFF;
            12'd   7: out = 16'hFFFF;
            12'd   8: out = 16'hFFFF;
            12'd   9: out = 16'hFFFF;
            12'd  10: out = 16'hFFFF;
            12'd  11: out = 16'hFFFF;
            12'd  12: out = 16'hFFFF;
            12'd  13: out = 16'hFFFF;
            12'd  14: out = 16'hFFFF;
            12'd  15: out = 16'hFFFF;
            12'd  16: out = 16'hFFFF;
            12'd  17: out = 16'hFFFF;
            12'd  18: out = 16'hFFFF;
            12'd  19: out = 16'hFFFF;
            12'd  20: out = 16'hFFFF;
            12'd  21: out = 16'hFFFF;
            12'd  22: out = 16'hFFFF;
            12'd  23: out = 16'hFFFF;
            12'd  24: out = 16'hFFFF;
            12'd  25: out = 16'hFFFF;
            12'd  26: out = 16'hFFFF;
            12'd  27: out = 16'hFFFF;
            12'd  28: out = 16'hFFFF;
            12'd  29: out = 16'hFFFF;
            12'd  30: out = 16'hFFFF;
            12'd  31: out = 16'hFFFF;
            12'd  32: out = 16'hFFFF;
            12'd  33: out = 16'hFFFF;
            12'd  34: out = 16'hFFFF;
            12'd  35: out = 16'hFFFF;
            12'd  36: out = 16'hFFFF;
            12'd  37: out = 16'hFFFF;
            12'd  38: out = 16'hFFFF;
            12'd  39: out = 16'hFFFF;
            12'd  40: out = 16'hFFFF;
            12'd  41: out = 16'hFFFF;
            12'd  42: out = 16'hFFFF;
            12'd  43: out = 16'hFFFF;
            12'd  44: out = 16'hFFFF;
            12'd  45: out = 16'hFFFF;
            12'd  46: out = 16'hFFFF;
            12'd  47: out = 16'hFFFF;
            12'd  48: out = 16'hFFFF;
            12'd  49: out = 16'hFFFF;
            12'd  50: out = 16'hFFFF;
            12'd  51: out = 16'hFFFF;
            12'd  52: out = 16'hFFFF;
            12'd  53: out = 16'hFFFF;
            12'd  54: out = 16'hFFFF;
            12'd  55: out = 16'hFFFF;
            12'd  56: out = 16'hFFFF;
            12'd  57: out = 16'hFFFF;
            12'd  58: out = 16'hFFFF;
            12'd  59: out = 16'hFFFF;
            12'd  60: out = 16'hFFFF;
            12'd  61: out = 16'hFFFF;
            12'd  62: out = 16'hFFFF;
            12'd  63: out = 16'hFFFF;
            12'd  64: out = 16'hFFFF;
            12'd  65: out = 16'hFFFF;
            12'd  66: out = 16'hFFFF;
            12'd  67: out = 16'hFFFF;
            12'd  68: out = 16'hFFFF;
            12'd  69: out = 16'hFFFF;
            12'd  70: out = 16'hFFFF;
            12'd  71: out = 16'hFFFF;
            12'd  72: out = 16'hFFFF;
            12'd  73: out = 16'hFFFF;
            12'd  74: out = 16'hFFFF;
            12'd  75: out = 16'hFFFF;
            12'd  76: out = 16'hFFFF;
            12'd  77: out = 16'hFFFF;
            12'd  78: out = 16'hFFFF;
            12'd  79: out = 16'hFFFF;
            12'd  80: out = 16'hFFFF;
            12'd  81: out = 16'hFFFF;
            12'd  82: out = 16'hFFFF;
            12'd  83: out = 16'hFFFF;
            12'd  84: out = 16'hFFFF;
            12'd  85: out = 16'hFFFF;
            12'd  86: out = 16'hFFFF;
            12'd  87: out = 16'hFFFF;
            12'd  88: out = 16'hFFFF;
            12'd  89: out = 16'hFFFF;
            12'd  90: out = 16'hFFFF;
            12'd  91: out = 16'hFFFF;
            12'd  92: out = 16'hFFFF;
            12'd  93: out = 16'hFFFF;
            12'd  94: out = 16'hFFFF;
            12'd  95: out = 16'hFFFF;
            12'd  96: out = 16'hFFFF;
            12'd  97: out = 16'hFFFF;
            12'd  98: out = 16'hFFFF;
            12'd  99: out = 16'hFFFF;
            12'd 100: out = 16'hFFFF;
            12'd 101: out = 16'hFFFF;
            12'd 102: out = 16'hFFFF;
            12'd 103: out = 16'hFFFF;
            12'd 104: out = 16'hFFFF;
            12'd 105: out = 16'hFFFF;
            12'd 106: out = 16'hFFFF;
            12'd 107: out = 16'hFFFF;
            12'd 108: out = 16'hFFFF;
            12'd 109: out = 16'hFFFF;
            12'd 110: out = 16'hFFFF;
            12'd 111: out = 16'hFFFF;
            12'd 112: out = 16'hFFFF;
            12'd 113: out = 16'hFFFF;
            12'd 114: out = 16'hFFFF;
            12'd 115: out = 16'hFFFF;
            12'd 116: out = 16'hFFFF;
            12'd 117: out = 16'hFFFF;
            12'd 118: out = 16'hFFFF;
            12'd 119: out = 16'hFFFF;
            12'd 120: out = 16'hFFFF;
            12'd 121: out = 16'hFFFF;
            12'd 122: out = 16'hFFFF;
            12'd 123: out = 16'hFFFF;
            12'd 124: out = 16'hFFFF;
            12'd 125: out = 16'hFFFF;
            12'd 126: out = 16'hFFFF;
            12'd 127: out = 16'hFFFF;
            12'd 128: out = 16'hFFFF;
            12'd 129: out = 16'hFFFF;
            12'd 130: out = 16'hFFFF;
            12'd 131: out = 16'hFFFF;
            12'd 132: out = 16'hFFFF;
            12'd 133: out = 16'hFFFF;
            12'd 134: out = 16'hFFFF;
            12'd 135: out = 16'hFFFF;
            12'd 136: out = 16'hFFFF;
            12'd 137: out = 16'hFFFF;
            12'd 138: out = 16'hFFFF;
            12'd 139: out = 16'hFFFF;
            12'd 140: out = 16'hFFFF;
            12'd 141: out = 16'hFFFF;
            12'd 142: out = 16'hFFFF;
            12'd 143: out = 16'hFFFF;
            12'd 144: out = 16'hFFFF;
            12'd 145: out = 16'hFFFF;
            12'd 146: out = 16'hFFFF;
            12'd 147: out = 16'hFFFF;
            12'd 148: out = 16'hFFFF;
            12'd 149: out = 16'hFFFF;
            12'd 150: out = 16'hFFFF;
            12'd 151: out = 16'hFFFF;
            12'd 152: out = 16'hFFFF;
            12'd 153: out = 16'hFFFF;
            12'd 154: out = 16'hFFFF;
            12'd 155: out = 16'hFFFF;
            12'd 156: out = 16'hFFFF;
            12'd 157: out = 16'hFFFF;
            12'd 158: out = 16'hFFFF;
            12'd 159: out = 16'hFFFF;
            12'd 160: out = 16'hFFFF;
            12'd 161: out = 16'hFFFF;
            12'd 162: out = 16'hFFFF;
            12'd 163: out = 16'hFFFF;
            12'd 164: out = 16'hFFFF;
            12'd 165: out = 16'hFFFF;
            12'd 166: out = 16'hFFFF;
            12'd 167: out = 16'hFFFF;
            12'd 168: out = 16'hFFFF;
            12'd 169: out = 16'hFFFF;
            12'd 170: out = 16'hFFFF;
            12'd 171: out = 16'hFFFF;
            12'd 172: out = 16'hFFFF;
            12'd 173: out = 16'hFFFF;
            12'd 174: out = 16'hFFFF;
            12'd 175: out = 16'hFFFF;
            12'd 176: out = 16'hFFFF;
            12'd 177: out = 16'hFFFF;
            12'd 178: out = 16'hFFFF;
            12'd 179: out = 16'hFFFF;
            12'd 180: out = 16'hFFFF;
            12'd 181: out = 16'hFFFF;
            12'd 182: out = 16'hFFFF;
            12'd 183: out = 16'hFFFF;
            12'd 184: out = 16'hFFFF;
            12'd 185: out = 16'hFFFF;
            12'd 186: out = 16'hFFFF;
            12'd 187: out = 16'hFFFF;
            12'd 188: out = 16'hFFFF;
            12'd 189: out = 16'hFFFF;
            12'd 190: out = 16'hFFFF;
            12'd 191: out = 16'hFFFF;
            12'd 192: out = 16'hFFFF;
            12'd 193: out = 16'hFFFF;
            12'd 194: out = 16'hFFFF;
            12'd 195: out = 16'hFFFF;
            12'd 196: out = 16'hFFFF;
            12'd 197: out = 16'hFFFF;
            12'd 198: out = 16'hFFFF;
            12'd 199: out = 16'hFFFF;
            12'd 200: out = 16'hFFFF;
            12'd 201: out = 16'hFFFF;
            12'd 202: out = 16'hFFFF;
            12'd 203: out = 16'hFFFF;
            12'd 204: out = 16'hFFFF;
            12'd 205: out = 16'hFFFF;
            12'd 206: out = 16'hFFFF;
            12'd 207: out = 16'hFFFF;
            12'd 208: out = 16'hFFFF;
            12'd 209: out = 16'hFFFF;
            12'd 210: out = 16'hFFFF;
            12'd 211: out = 16'hFFFF;
            12'd 212: out = 16'hFFFF;
            12'd 213: out = 16'hFFFF;
            12'd 214: out = 16'hFFFF;
            12'd 215: out = 16'hFFFF;
            12'd 216: out = 16'hFFFF;
            12'd 217: out = 16'hFFFF;
            12'd 218: out = 16'hFFFF;
            12'd 219: out = 16'hFFFF;
            12'd 220: out = 16'hFFFF;
            12'd 221: out = 16'hFFFF;
            12'd 222: out = 16'hFFFF;
            12'd 223: out = 16'hFFFF;
            12'd 224: out = 16'hFFFF;
            12'd 225: out = 16'hFFFF;
            12'd 226: out = 16'hFFFF;
            12'd 227: out = 16'hFFFF;
            12'd 228: out = 16'hFFFF;
            12'd 229: out = 16'hFFFF;
            12'd 230: out = 16'hFFFF;
            12'd 231: out = 16'hFFFF;
            12'd 232: out = 16'hFFFF;
            12'd 233: out = 16'hFFFF;
            12'd 234: out = 16'hFFFF;
            12'd 235: out = 16'hFFFF;
            12'd 236: out = 16'hFFFF;
            12'd 237: out = 16'hFFFF;
            12'd 238: out = 16'hFFFF;
            12'd 239: out = 16'hFFFF;
            12'd 240: out = 16'hFFFF;
            12'd 241: out = 16'hFFFF;
            12'd 242: out = 16'hFFFF;
            12'd 243: out = 16'hFFFF;
            12'd 244: out = 16'hFFFF;
            12'd 245: out = 16'hFFFF;
            12'd 246: out = 16'hFFFF;
            12'd 247: out = 16'hFFFF;
            12'd 248: out = 16'hFFFF;
            12'd 249: out = 16'hFFFF;
            12'd 250: out = 16'hFFFF;
            12'd 251: out = 16'hFFFF;
            12'd 252: out = 16'hFFFF;
            12'd 253: out = 16'hFFFF;
            12'd 254: out = 16'hFFFF;
            12'd 255: out = 16'hFFFF;
            12'd 256: out = 16'hFFFF;
            12'd 257: out = 16'hFFFF;
            12'd 258: out = 16'hFFFF;
            12'd 259: out = 16'hFFFF;
            12'd 260: out = 16'hFFFF;
            12'd 261: out = 16'hFFFF;
            12'd 262: out = 16'hFFFF;
            12'd 263: out = 16'hFFFF;
            12'd 264: out = 16'hFFFF;
            12'd 265: out = 16'hFFFF;
            12'd 266: out = 16'hFFFF;
            12'd 267: out = 16'hFFFF;
            12'd 268: out = 16'hFFFF;
            12'd 269: out = 16'hFFFF;
            12'd 270: out = 16'hFFFF;
            12'd 271: out = 16'hFFFF;
            12'd 272: out = 16'hFFFF;
            12'd 273: out = 16'hFFFF;
            12'd 274: out = 16'hFFFF;
            12'd 275: out = 16'hFFFF;
            12'd 276: out = 16'hFFFF;
            12'd 277: out = 16'hFFFF;
            12'd 278: out = 16'hFFFF;
            12'd 279: out = 16'hFFFF;
            12'd 280: out = 16'hFFFF;
            12'd 281: out = 16'hFFFF;
            12'd 282: out = 16'hFFFF;
            12'd 283: out = 16'hFFFF;
            12'd 284: out = 16'hFFFF;
            12'd 285: out = 16'hFFFF;
            12'd 286: out = 16'hFFFF;
            12'd 287: out = 16'hFFFF;
            12'd 288: out = 16'hFFFF;
            12'd 289: out = 16'hFFFF;
            12'd 290: out = 16'hFFFF;
            12'd 291: out = 16'hFFFF;
            12'd 292: out = 16'hFFFF;
            12'd 293: out = 16'hFFFF;
            12'd 294: out = 16'hFFFF;
            12'd 295: out = 16'hFFFF;
            12'd 296: out = 16'hFFFF;
            12'd 297: out = 16'hFFFF;
            12'd 298: out = 16'hFFFF;
            12'd 299: out = 16'hFFFF;
            12'd 300: out = 16'hFFFF;
            12'd 301: out = 16'hFFFF;
            12'd 302: out = 16'hFFFF;
            12'd 303: out = 16'hFFFF;
            12'd 304: out = 16'hFFFF;
            12'd 305: out = 16'hFFFF;
            12'd 306: out = 16'hFFFF;
            12'd 307: out = 16'hFFFF;
            12'd 308: out = 16'hFFFF;
            12'd 309: out = 16'hFFFF;
            12'd 310: out = 16'hFFFF;
            12'd 311: out = 16'hFFFF;
            12'd 312: out = 16'hFFFF;
            12'd 313: out = 16'hFFFF;
            12'd 314: out = 16'hFFFF;
            12'd 315: out = 16'hFFFF;
            12'd 316: out = 16'hFFFF;
            12'd 317: out = 16'hFFFF;
            12'd 318: out = 16'hFFFF;
            12'd 319: out = 16'hFFFF;
            12'd 320: out = 16'hFFFF;
            12'd 321: out = 16'hFFFF;
            12'd 322: out = 16'hFFFF;
            12'd 323: out = 16'hFFFF;
            12'd 324: out = 16'hFFFF;
            12'd 325: out = 16'hFFFF;
            12'd 326: out = 16'hFFFF;
            12'd 327: out = 16'hFFFF;
            12'd 328: out = 16'hFFFF;
            12'd 329: out = 16'hFFFF;
            12'd 330: out = 16'hFFFF;
            12'd 331: out = 16'hFFFF;
            12'd 332: out = 16'hFFFF;
            12'd 333: out = 16'hFFFF;
            12'd 334: out = 16'hFFFF;
            12'd 335: out = 16'hFFFF;
            12'd 336: out = 16'hFFFF;
            12'd 337: out = 16'hFFFF;
            12'd 338: out = 16'hFFFF;
            12'd 339: out = 16'hFFFF;
            12'd 340: out = 16'hFFFF;
            12'd 341: out = 16'hFFFF;
            12'd 342: out = 16'hFFFF;
            12'd 343: out = 16'hFFFF;
            12'd 344: out = 16'hFFFF;
            12'd 345: out = 16'hFFFF;
            12'd 346: out = 16'hFFFF;
            12'd 347: out = 16'hFFFF;
            12'd 348: out = 16'hFFFF;
            12'd 349: out = 16'hFFFF;
            12'd 350: out = 16'hFFFF;
            12'd 351: out = 16'hFFFF;
            12'd 352: out = 16'hFFFF;
            12'd 353: out = 16'hFFFF;
            12'd 354: out = 16'hFFFF;
            12'd 355: out = 16'hFFFF;
            12'd 356: out = 16'hFFFF;
            12'd 357: out = 16'hFFFF;
            12'd 358: out = 16'hFFFF;
            12'd 359: out = 16'hFFFF;
            12'd 360: out = 16'hFFFF;
            12'd 361: out = 16'hFFFF;
            12'd 362: out = 16'hFFFF;
            12'd 363: out = 16'hFFFF;
            12'd 364: out = 16'hFFFF;
            12'd 365: out = 16'hFFFF;
            12'd 366: out = 16'hFFFF;
            12'd 367: out = 16'hFFFF;
            12'd 368: out = 16'hFFFF;
            12'd 369: out = 16'hFFFF;
            12'd 370: out = 16'hFFFF;
            12'd 371: out = 16'hFFFF;
            12'd 372: out = 16'hFFFF;
            12'd 373: out = 16'hFFFF;
            12'd 374: out = 16'hFFFF;
            12'd 375: out = 16'hFFFF;
            12'd 376: out = 16'hFFFF;
            12'd 377: out = 16'hFFFF;
            12'd 378: out = 16'hFFFF;
            12'd 379: out = 16'hFFFF;
            12'd 380: out = 16'hFFFF;
            12'd 381: out = 16'hFFFF;
            12'd 382: out = 16'hFFFF;
            12'd 383: out = 16'hFFFF;
            12'd 384: out = 16'hFFFF;
            12'd 385: out = 16'hFFFF;
            12'd 386: out = 16'hFFFF;
            12'd 387: out = 16'hFFFF;
            12'd 388: out = 16'hFFFF;
            12'd 389: out = 16'hFFFF;
            12'd 390: out = 16'hFFFF;
            12'd 391: out = 16'hFFFF;
            12'd 392: out = 16'hFFFF;
            12'd 393: out = 16'hFFFF;
            12'd 394: out = 16'hFFFF;
            12'd 395: out = 16'hFFFF;
            12'd 396: out = 16'hFFFF;
            12'd 397: out = 16'hFFFF;
            12'd 398: out = 16'hFFFF;
            12'd 399: out = 16'hFFFF;
            12'd 400: out = 16'hFFFF;
            12'd 401: out = 16'hFFFF;
            12'd 402: out = 16'hFFFF;
            12'd 403: out = 16'hFFFF;
            12'd 404: out = 16'hFFFF;
            12'd 405: out = 16'hFFFF;
            12'd 406: out = 16'hFFFF;
            12'd 407: out = 16'hFFFF;
            12'd 408: out = 16'hFFFF;
            12'd 409: out = 16'hFFFF;
            12'd 410: out = 16'hFFFF;
            12'd 411: out = 16'hFFFF;
            12'd 412: out = 16'hFFFF;
            12'd 413: out = 16'hFFFF;
            12'd 414: out = 16'hFFFF;
            12'd 415: out = 16'hFFFF;
            12'd 416: out = 16'hFFFF;
            12'd 417: out = 16'hFFFF;
            12'd 418: out = 16'hFFFF;
            12'd 419: out = 16'hFFFF;
            12'd 420: out = 16'hFFFF;
            12'd 421: out = 16'hFFFF;
            12'd 422: out = 16'hFFFF;
            12'd 423: out = 16'hFFFF;
            12'd 424: out = 16'hFFFF;
            12'd 425: out = 16'hFFFF;
            12'd 426: out = 16'hFFFF;
            12'd 427: out = 16'hFFFF;
            12'd 428: out = 16'hFFFF;
            12'd 429: out = 16'hFFFF;
            12'd 430: out = 16'hFFFF;
            12'd 431: out = 16'hFFFF;
            12'd 432: out = 16'hFFFF;
            12'd 433: out = 16'hFFFF;
            12'd 434: out = 16'hFFFF;
            12'd 435: out = 16'hFFFF;
            12'd 436: out = 16'hFFFF;
            12'd 437: out = 16'hFFFF;
            12'd 438: out = 16'hFFFF;
            12'd 439: out = 16'hFFFF;
            12'd 440: out = 16'hFFFF;
            12'd 441: out = 16'hFFFF;
            12'd 442: out = 16'hFFFF;
            12'd 443: out = 16'hFFFF;
            12'd 444: out = 16'hFFFF;
            12'd 445: out = 16'hFFFF;
            12'd 446: out = 16'hFFFF;
            12'd 447: out = 16'hFFFF;
            12'd 448: out = 16'hFFFF;
            12'd 449: out = 16'hFFFF;
            12'd 450: out = 16'hFFFF;
            12'd 451: out = 16'hFFFF;
            12'd 452: out = 16'hFFFF;
            12'd 453: out = 16'hFFFF;
            12'd 454: out = 16'hFFFF;
            12'd 455: out = 16'hFFFF;
            12'd 456: out = 16'hFFFF;
            12'd 457: out = 16'hFFFF;
            12'd 458: out = 16'hFFFF;
            12'd 459: out = 16'hFFFF;
            12'd 460: out = 16'hFFFF;
            12'd 461: out = 16'hFFFF;
            12'd 462: out = 16'hFFFF;
            12'd 463: out = 16'hFFFF;
            12'd 464: out = 16'hFFFF;
            12'd 465: out = 16'hFFFF;
            12'd 466: out = 16'hFFFF;
            12'd 467: out = 16'hFFFF;
            12'd 468: out = 16'hFFFF;
            12'd 469: out = 16'hFFFF;
            12'd 470: out = 16'hFFFF;
            12'd 471: out = 16'hFFFF;
            12'd 472: out = 16'hFFFF;
            12'd 473: out = 16'hFFFF;
            12'd 474: out = 16'hFFFF;
            12'd 475: out = 16'hFFFF;
            12'd 476: out = 16'hFFFF;
            12'd 477: out = 16'hFFFF;
            12'd 478: out = 16'hFFFF;
            12'd 479: out = 16'hFFFF;
            12'd 480: out = 16'hFFFF;
            12'd 481: out = 16'hFFFF;
            12'd 482: out = 16'hFFFF;
            12'd 483: out = 16'hFFFF;
            12'd 484: out = 16'hFFFF;
            12'd 485: out = 16'hFFFF;
            12'd 486: out = 16'hFFFF;
            12'd 487: out = 16'hFFFF;
            12'd 488: out = 16'hFFFF;
            12'd 489: out = 16'hFFFF;
            12'd 490: out = 16'hFFFF;
            12'd 491: out = 16'hFFFF;
            12'd 492: out = 16'hFFFF;
            12'd 493: out = 16'hFFFF;
            12'd 494: out = 16'hFFFF;
            12'd 495: out = 16'hFFFF;
            12'd 496: out = 16'hFFFF;
            12'd 497: out = 16'hFFFF;
            12'd 498: out = 16'hFFFF;
            12'd 499: out = 16'hFFFF;
            12'd 500: out = 16'hFFFF;
            12'd 501: out = 16'hFFFF;
            12'd 502: out = 16'hFFFF;
            12'd 503: out = 16'hFFFF;
            12'd 504: out = 16'hFFFF;
            12'd 505: out = 16'hFFFF;
            12'd 506: out = 16'hFFFF;
            12'd 507: out = 16'hFFFF;
            12'd 508: out = 16'hFFFF;
            12'd 509: out = 16'hFFFF;
            12'd 510: out = 16'hFFFF;
            12'd 511: out = 16'hFFFF;
            12'd 512: out = 16'hFFFF;
            12'd 513: out = 16'hFFFF;
            12'd 514: out = 16'hFFFF;
            12'd 515: out = 16'hFFFF;
            12'd 516: out = 16'hFFFF;
            12'd 517: out = 16'hFFFF;
            12'd 518: out = 16'hFFFF;
            12'd 519: out = 16'hFFFF;
            12'd 520: out = 16'hFFFF;
            12'd 521: out = 16'hFFFF;
            12'd 522: out = 16'hFFFF;
            12'd 523: out = 16'hFFFF;
            12'd 524: out = 16'hFFFF;
            12'd 525: out = 16'hFFFF;
            12'd 526: out = 16'hFFFF;
            12'd 527: out = 16'hFFFF;
            12'd 528: out = 16'hFFFF;
            12'd 529: out = 16'hFFFF;
            12'd 530: out = 16'hFFFF;
            12'd 531: out = 16'hFFFF;
            12'd 532: out = 16'hFFFF;
            12'd 533: out = 16'hFFFF;
            12'd 534: out = 16'hFFFF;
            12'd 535: out = 16'hFFFF;
            12'd 536: out = 16'hFFFF;
            12'd 537: out = 16'hFFFF;
            12'd 538: out = 16'hFFFF;
            12'd 539: out = 16'hFFFF;
            12'd 540: out = 16'hFFFF;
            12'd 541: out = 16'hFFFF;
            12'd 542: out = 16'hFFFF;
            12'd 543: out = 16'hFFFF;
            12'd 544: out = 16'hFFFF;
            12'd 545: out = 16'hFFFF;
            12'd 546: out = 16'hFFFF;
            12'd 547: out = 16'hFFFF;
            12'd 548: out = 16'hFFFF;
            12'd 549: out = 16'hFFFF;
            12'd 550: out = 16'hFFFF;
            12'd 551: out = 16'hFFFF;
            12'd 552: out = 16'hFFFF;
            12'd 553: out = 16'hFFFF;
            12'd 554: out = 16'hFFFF;
            12'd 555: out = 16'hFFFF;
            12'd 556: out = 16'hFFFF;
            12'd 557: out = 16'hFFFF;
            12'd 558: out = 16'hFFFF;
            12'd 559: out = 16'hFFFF;
            12'd 560: out = 16'hFFFF;
            12'd 561: out = 16'hFFFF;
            12'd 562: out = 16'hFFFF;
            12'd 563: out = 16'hFFFF;
            12'd 564: out = 16'hFFFF;
            12'd 565: out = 16'hFFFF;
            12'd 566: out = 16'hFFFF;
            12'd 567: out = 16'hFFFF;
            12'd 568: out = 16'hFFFF;
            12'd 569: out = 16'hFFFF;
            12'd 570: out = 16'hFFFF;
            12'd 571: out = 16'hFFFF;
            12'd 572: out = 16'hFFFF;
            12'd 573: out = 16'hFFFF;
            12'd 574: out = 16'hFFFF;
            12'd 575: out = 16'hFFFF;
            12'd 576: out = 16'hFFFF;
            12'd 577: out = 16'hFFFF;
            12'd 578: out = 16'hFFFF;
            12'd 579: out = 16'hFFFF;
            12'd 580: out = 16'hFFFF;
            12'd 581: out = 16'hFFFF;
            12'd 582: out = 16'hFFFF;
            12'd 583: out = 16'hFFFF;
            12'd 584: out = 16'hFFFF;
            12'd 585: out = 16'hFFFF;
            12'd 586: out = 16'hFFFF;
            12'd 587: out = 16'hFFFF;
            12'd 588: out = 16'hFFFF;
            12'd 589: out = 16'hFFFF;
            12'd 590: out = 16'hFFFF;
            12'd 591: out = 16'hFFFF;
            12'd 592: out = 16'hFFFF;
            12'd 593: out = 16'hFFFF;
            12'd 594: out = 16'hFFFF;
            12'd 595: out = 16'hFFFF;
            12'd 596: out = 16'hFFFF;
            12'd 597: out = 16'hFFFF;
            12'd 598: out = 16'hFFFF;
            12'd 599: out = 16'hFFFF;
            12'd 600: out = 16'hFFFF;
            12'd 601: out = 16'hFFFF;
            12'd 602: out = 16'hFFFF;
            12'd 603: out = 16'hFFFF;
            12'd 604: out = 16'hFFFF;
            12'd 605: out = 16'hFFFF;
            12'd 606: out = 16'hFFFF;
            12'd 607: out = 16'hFFFF;
            12'd 608: out = 16'hFFFF;
            12'd 609: out = 16'hFFFF;
            12'd 610: out = 16'hFFFF;
            12'd 611: out = 16'hFFFF;
            12'd 612: out = 16'hFFFF;
            12'd 613: out = 16'hFFFF;
            12'd 614: out = 16'hFFFF;
            12'd 615: out = 16'hFFFF;
            12'd 616: out = 16'hFFFF;
            12'd 617: out = 16'hFFFF;
            12'd 618: out = 16'hFFFF;
            12'd 619: out = 16'hFFFF;
            12'd 620: out = 16'hFFFF;
            12'd 621: out = 16'hFFFF;
            12'd 622: out = 16'hFFFF;
            12'd 623: out = 16'hFFFF;
            12'd 624: out = 16'hFFFF;
            12'd 625: out = 16'hFFFF;
            12'd 626: out = 16'hFFFF;
            12'd 627: out = 16'hFFFF;
            12'd 628: out = 16'hFFFF;
            12'd 629: out = 16'hFFFF;
            12'd 630: out = 16'hFFFF;
            12'd 631: out = 16'hFFFF;
            12'd 632: out = 16'hFFFF;
            12'd 633: out = 16'hFFFF;
            12'd 634: out = 16'hFFFF;
            12'd 635: out = 16'hFFFF;
            12'd 636: out = 16'hFFFF;
            12'd 637: out = 16'hFFFF;
            12'd 638: out = 16'hFFFF;
            12'd 639: out = 16'hFFFF;
            12'd 640: out = 16'hFFFF;
            12'd 641: out = 16'hFFFF;
            12'd 642: out = 16'hFFFF;
            12'd 643: out = 16'hFFFF;
            12'd 644: out = 16'hFFFF;
            12'd 645: out = 16'hFFFF;
            12'd 646: out = 16'hFFFF;
            12'd 647: out = 16'hFFFF;
            12'd 648: out = 16'hFFFF;
            12'd 649: out = 16'hFFFF;
            12'd 650: out = 16'hFFFF;
            12'd 651: out = 16'hFFFF;
            12'd 652: out = 16'hFFFF;
            12'd 653: out = 16'hFFFF;
            12'd 654: out = 16'hFFFF;
            12'd 655: out = 16'hFFFF;
            12'd 656: out = 16'hFFFF;
            12'd 657: out = 16'hFFFF;
            12'd 658: out = 16'hFFFF;
            12'd 659: out = 16'hFFFF;
            12'd 660: out = 16'hFFFF;
            12'd 661: out = 16'hFFFF;
            12'd 662: out = 16'hFFFF;
            12'd 663: out = 16'hFFFF;
            12'd 664: out = 16'hFFFF;
            12'd 665: out = 16'hFFFF;
            12'd 666: out = 16'hFFFF;
            12'd 667: out = 16'hFFFF;
            12'd 668: out = 16'hFFFF;
            12'd 669: out = 16'hFFFF;
            12'd 670: out = 16'hFFFF;
            12'd 671: out = 16'hFFFF;
            12'd 672: out = 16'hFFFF;
            12'd 673: out = 16'hFFFF;
            12'd 674: out = 16'hFFFF;
            12'd 675: out = 16'hFFFF;
            12'd 676: out = 16'hFFFF;
            12'd 677: out = 16'hFFFF;
            12'd 678: out = 16'hFFFF;
            12'd 679: out = 16'hFFFF;
            12'd 680: out = 16'hFFFF;
            12'd 681: out = 16'hFFFF;
            12'd 682: out = 16'hFFFF;
            12'd 683: out = 16'hFFFF;
            12'd 684: out = 16'hFFFF;
            12'd 685: out = 16'hFFFF;
            12'd 686: out = 16'hFFFF;
            12'd 687: out = 16'hFFFF;
            12'd 688: out = 16'hFFFF;
            12'd 689: out = 16'hFFFF;
            12'd 690: out = 16'hFFFF;
            12'd 691: out = 16'hFFFF;
            12'd 692: out = 16'hFFFF;
            12'd 693: out = 16'hFFFF;
            12'd 694: out = 16'hFFFF;
            12'd 695: out = 16'hFFFF;
            12'd 696: out = 16'hFFFF;
            12'd 697: out = 16'hFFFF;
            12'd 698: out = 16'hFFFF;
            12'd 699: out = 16'hFFFF;
            12'd 700: out = 16'hFFFF;
            12'd 701: out = 16'hFFFF;
            12'd 702: out = 16'hFFFF;
            12'd 703: out = 16'hFFFF;
            12'd 704: out = 16'hFFFF;
            12'd 705: out = 16'hFFFF;
            12'd 706: out = 16'hFFFF;
            12'd 707: out = 16'hFFFF;
            12'd 708: out = 16'hFFFF;
            12'd 709: out = 16'hFFFF;
            12'd 710: out = 16'hFFFF;
            12'd 711: out = 16'hFFFF;
            12'd 712: out = 16'hFFFF;
            12'd 713: out = 16'hFFFF;
            12'd 714: out = 16'hFFFF;
            12'd 715: out = 16'hFFFF;
            12'd 716: out = 16'hFFFF;
            12'd 717: out = 16'hFFFF;
            12'd 718: out = 16'hFFFF;
            12'd 719: out = 16'hFFFF;
            12'd 720: out = 16'hFFFF;
            12'd 721: out = 16'hFFFF;
            12'd 722: out = 16'hFFFF;
            12'd 723: out = 16'hFFFF;
            12'd 724: out = 16'hFFFF;
            12'd 725: out = 16'hFFFF;
            12'd 726: out = 16'hFFFF;
            12'd 727: out = 16'hFFFF;
            12'd 728: out = 16'hFFFF;
            12'd 729: out = 16'hFFFF;
            12'd 730: out = 16'hFFFF;
            12'd 731: out = 16'hFFFF;
            12'd 732: out = 16'hFFFF;
            12'd 733: out = 16'hFFFF;
            12'd 734: out = 16'hFFFF;
            12'd 735: out = 16'hFFFF;
            12'd 736: out = 16'hFFFF;
            12'd 737: out = 16'hFFFF;
            12'd 738: out = 16'hFFFF;
            12'd 739: out = 16'hFFFF;
            12'd 740: out = 16'hFFFF;
            12'd 741: out = 16'hFFFF;
            12'd 742: out = 16'hFFFF;
            12'd 743: out = 16'hFFFF;
            12'd 744: out = 16'hFFFF;
            12'd 745: out = 16'hFFFF;
            12'd 746: out = 16'hFFFF;
            12'd 747: out = 16'hFFFF;
            12'd 748: out = 16'hFFFF;
            12'd 749: out = 16'hFFFF;
            12'd 750: out = 16'hFFFF;
            12'd 751: out = 16'hFFFF;
            12'd 752: out = 16'hFFFF;
            12'd 753: out = 16'hFFFF;
            12'd 754: out = 16'hFFFF;
            12'd 755: out = 16'hFFFF;
            12'd 756: out = 16'hFFFF;
            12'd 757: out = 16'hFFFF;
            12'd 758: out = 16'hFFFF;
            12'd 759: out = 16'hFFFF;
            12'd 760: out = 16'hFFFF;
            12'd 761: out = 16'hFFFF;
            12'd 762: out = 16'hFFFF;
            12'd 763: out = 16'hFFFF;
            12'd 764: out = 16'hFFFF;
            12'd 765: out = 16'hFFFF;
            12'd 766: out = 16'hFFFF;
            12'd 767: out = 16'hFFFF;
            12'd 768: out = 16'hFFFF;
            12'd 769: out = 16'hFFFF;
            12'd 770: out = 16'hFFFF;
            12'd 771: out = 16'hFFFF;
            12'd 772: out = 16'hFFFF;
            12'd 773: out = 16'hFFFF;
            12'd 774: out = 16'hFFFF;
            12'd 775: out = 16'hFFFF;
            12'd 776: out = 16'hFFFF;
            12'd 777: out = 16'hFFFF;
            12'd 778: out = 16'hFFFF;
            12'd 779: out = 16'hFFFF;
            12'd 780: out = 16'hFFFF;
            12'd 781: out = 16'hFFFF;
            12'd 782: out = 16'hFFFF;
            12'd 783: out = 16'hFFFF;
            12'd 784: out = 16'hFFFF;
            12'd 785: out = 16'hFFFF;
            12'd 786: out = 16'hFFFF;
            12'd 787: out = 16'hFFFF;
            12'd 788: out = 16'hFFFF;
            12'd 789: out = 16'hFFFF;
            12'd 790: out = 16'hFFFF;
            12'd 791: out = 16'hFFFF;
            12'd 792: out = 16'hFFFF;
            12'd 793: out = 16'hFFFF;
            12'd 794: out = 16'hFFFF;
            12'd 795: out = 16'hFFFF;
            12'd 796: out = 16'hFFFF;
            12'd 797: out = 16'hFFFF;
            12'd 798: out = 16'hFFFF;
            12'd 799: out = 16'hFFFF;
            12'd 800: out = 16'hFFFF;
            12'd 801: out = 16'hFFFF;
            12'd 802: out = 16'hFFFF;
            12'd 803: out = 16'hFFFF;
            12'd 804: out = 16'hFFFF;
            12'd 805: out = 16'hFFFF;
            12'd 806: out = 16'hFFFF;
            12'd 807: out = 16'hFFFF;
            12'd 808: out = 16'hFFFF;
            12'd 809: out = 16'hFFFF;
            12'd 810: out = 16'hFFFF;
            12'd 811: out = 16'hFFFF;
            12'd 812: out = 16'hFFFF;
            12'd 813: out = 16'hFFFF;
            12'd 814: out = 16'hFFFF;
            12'd 815: out = 16'hFFFF;
            12'd 816: out = 16'hFFFF;
            12'd 817: out = 16'hFFFF;
            12'd 818: out = 16'hFFFF;
            12'd 819: out = 16'hFFFF;
            12'd 820: out = 16'hFFFF;
            12'd 821: out = 16'hFFFF;
            12'd 822: out = 16'hFFFF;
            12'd 823: out = 16'hFFFF;
            12'd 824: out = 16'hFFFF;
            12'd 825: out = 16'hFFFF;
            12'd 826: out = 16'hFFFF;
            12'd 827: out = 16'hFFFF;
            12'd 828: out = 16'hFFFF;
            12'd 829: out = 16'hFFFF;
            12'd 830: out = 16'hFFFF;
            12'd 831: out = 16'hFFFF;
            12'd 832: out = 16'hFFFF;
            12'd 833: out = 16'hFFFF;
            12'd 834: out = 16'hFFFF;
            12'd 835: out = 16'hFFFF;
            12'd 836: out = 16'hFFFF;
            12'd 837: out = 16'hFFFF;
            12'd 838: out = 16'hFFFF;
            12'd 839: out = 16'hFFFF;
            12'd 840: out = 16'hFFFF;
            12'd 841: out = 16'hFFFF;
            12'd 842: out = 16'hFFFF;
            12'd 843: out = 16'hFFFF;
            12'd 844: out = 16'hFFFF;
            12'd 845: out = 16'hFFFF;
            12'd 846: out = 16'hFFFF;
            12'd 847: out = 16'hFFFF;
            12'd 848: out = 16'hFFFF;
            12'd 849: out = 16'hFFFF;
            12'd 850: out = 16'hFFFF;
            12'd 851: out = 16'hFFFF;
            12'd 852: out = 16'hFFFF;
            12'd 853: out = 16'hFFFF;
            12'd 854: out = 16'hFFFF;
            12'd 855: out = 16'hFFFF;
            12'd 856: out = 16'hFFFF;
            12'd 857: out = 16'hFFFF;
            12'd 858: out = 16'hFFFF;
            12'd 859: out = 16'hFFFF;
            12'd 860: out = 16'hFFFF;
            12'd 861: out = 16'hFFFF;
            12'd 862: out = 16'hFFFF;
            12'd 863: out = 16'hFFFF;
            12'd 864: out = 16'hFFFF;
            12'd 865: out = 16'hFFFF;
            12'd 866: out = 16'hFFFF;
            12'd 867: out = 16'hFFFF;
            12'd 868: out = 16'hFFFF;
            12'd 869: out = 16'hFFFF;
            12'd 870: out = 16'hFFFF;
            12'd 871: out = 16'hFFFF;
            12'd 872: out = 16'hFFFF;
            12'd 873: out = 16'hFFFF;
            12'd 874: out = 16'hFFFF;
            12'd 875: out = 16'hFFFF;
            12'd 876: out = 16'hFFFF;
            12'd 877: out = 16'hFFFF;
            12'd 878: out = 16'hFFFF;
            12'd 879: out = 16'hFFFF;
            12'd 880: out = 16'hFFFF;
            12'd 881: out = 16'hFFFF;
            12'd 882: out = 16'hFFFF;
            12'd 883: out = 16'hFFFF;
            12'd 884: out = 16'hFFFF;
            12'd 885: out = 16'hFFFF;
            12'd 886: out = 16'hFFFF;
            12'd 887: out = 16'hFFFF;
            12'd 888: out = 16'hFFFF;
            12'd 889: out = 16'hFFFF;
            12'd 890: out = 16'hFFFF;
            12'd 891: out = 16'hFFFF;
            12'd 892: out = 16'hFFFF;
            12'd 893: out = 16'hFFFF;
            12'd 894: out = 16'hFFFF;
            12'd 895: out = 16'hFFFF;
            12'd 896: out = 16'hFFFF;
            12'd 897: out = 16'hFFFF;
            12'd 898: out = 16'hFFFF;
            12'd 899: out = 16'hFFFF;
            12'd 900: out = 16'hFFFF;
            12'd 901: out = 16'hFFFF;
            12'd 902: out = 16'hFFFF;
            12'd 903: out = 16'hFFFF;
            12'd 904: out = 16'hFFFF;
            12'd 905: out = 16'hFFFF;
            12'd 906: out = 16'hFFFF;
            12'd 907: out = 16'hFFFF;
            12'd 908: out = 16'hFFFF;
            12'd 909: out = 16'hFFFF;
            12'd 910: out = 16'hFFFF;
            12'd 911: out = 16'hFFFF;
            12'd 912: out = 16'hFFFF;
            12'd 913: out = 16'hFFFF;
            12'd 914: out = 16'hFFFF;
            12'd 915: out = 16'hFFFF;
            12'd 916: out = 16'hFFFF;
            12'd 917: out = 16'hFFFF;
            12'd 918: out = 16'hFFFF;
            12'd 919: out = 16'hFFFF;
            12'd 920: out = 16'hFFFF;
            12'd 921: out = 16'hFFFF;
            12'd 922: out = 16'hFFFF;
            12'd 923: out = 16'hFFFF;
            12'd 924: out = 16'hFFFF;
            12'd 925: out = 16'hFFFF;
            12'd 926: out = 16'hFFFF;
            12'd 927: out = 16'hFFFF;
            12'd 928: out = 16'hFFFF;
            12'd 929: out = 16'hFFFF;
            12'd 930: out = 16'hFFFF;
            12'd 931: out = 16'hFFFF;
            12'd 932: out = 16'hFFFF;
            12'd 933: out = 16'hFFFF;
            12'd 934: out = 16'hFFFF;
            12'd 935: out = 16'hFFFF;
            12'd 936: out = 16'hFFFF;
            12'd 937: out = 16'hFFFF;
            12'd 938: out = 16'hFFFF;
            12'd 939: out = 16'hFFFF;
            12'd 940: out = 16'hFFFF;
            12'd 941: out = 16'hFFFF;
            12'd 942: out = 16'hFFFF;
            12'd 943: out = 16'hFFFF;
            12'd 944: out = 16'hFFFF;
            12'd 945: out = 16'hFFFF;
            12'd 946: out = 16'hFFFF;
            12'd 947: out = 16'hFFFF;
            12'd 948: out = 16'hFFFF;
            12'd 949: out = 16'hFFFF;
            12'd 950: out = 16'hFFFF;
            12'd 951: out = 16'hFFFF;
            12'd 952: out = 16'hFFFF;
            12'd 953: out = 16'hFFFF;
            12'd 954: out = 16'hFFFF;
            12'd 955: out = 16'hFFFF;
            12'd 956: out = 16'hFFFF;
            12'd 957: out = 16'hFFFF;
            12'd 958: out = 16'hFFFF;
            12'd 959: out = 16'hFFFF;
            12'd 960: out = 16'hFFFF;
            12'd 961: out = 16'hFFFF;
            12'd 962: out = 16'hFFFF;
            12'd 963: out = 16'hFFFF;
            12'd 964: out = 16'hFFFF;
            12'd 965: out = 16'hFFFF;
            12'd 966: out = 16'hFFFF;
            12'd 967: out = 16'hFFFF;
            12'd 968: out = 16'hFFFF;
            12'd 969: out = 16'hFFFF;
            12'd 970: out = 16'hFFFF;
            12'd 971: out = 16'hFFFF;
            12'd 972: out = 16'hFFFF;
            12'd 973: out = 16'hFFFF;
            12'd 974: out = 16'hFFFF;
            12'd 975: out = 16'hFFFF;
            12'd 976: out = 16'hFFFF;
            12'd 977: out = 16'hFFFF;
            12'd 978: out = 16'hFFFF;
            12'd 979: out = 16'hFFFF;
            12'd 980: out = 16'hFFFF;
            12'd 981: out = 16'hFFFF;
            12'd 982: out = 16'hFFFF;
            12'd 983: out = 16'hFFFF;
            12'd 984: out = 16'hFFFF;
            12'd 985: out = 16'hFFFF;
            12'd 986: out = 16'hFFFF;
            12'd 987: out = 16'hFFFF;
            12'd 988: out = 16'hFFFF;
            12'd 989: out = 16'hFFFF;
            12'd 990: out = 16'hFFFF;
            12'd 991: out = 16'hFFFF;
            12'd 992: out = 16'hFFFF;
            12'd 993: out = 16'hFFFF;
            12'd 994: out = 16'hFFFF;
            12'd 995: out = 16'hFFFF;
            12'd 996: out = 16'hFFFF;
            12'd 997: out = 16'hFFFF;
            12'd 998: out = 16'hFFFF;
            12'd 999: out = 16'hFFFF;
            12'd1000: out = 16'hFFFF;
            12'd1001: out = 16'hFFFF;
            12'd1002: out = 16'hFFFF;
            12'd1003: out = 16'hFFFF;
            12'd1004: out = 16'hFFFF;
            12'd1005: out = 16'hFFFF;
            12'd1006: out = 16'hFFFF;
            12'd1007: out = 16'hFFFF;
            12'd1008: out = 16'hFFFF;
            12'd1009: out = 16'hFFFF;
            12'd1010: out = 16'hFFFF;
            12'd1011: out = 16'hFFFF;
            12'd1012: out = 16'hFFFF;
            12'd1013: out = 16'hFFFF;
            12'd1014: out = 16'hFFFF;
            12'd1015: out = 16'hFFFF;
            12'd1016: out = 16'hFFFF;
            12'd1017: out = 16'hFFFF;
            12'd1018: out = 16'hFFFF;
            12'd1019: out = 16'hFFFF;
            12'd1020: out = 16'hFFFF;
            12'd1021: out = 16'hFFFF;
            12'd1022: out = 16'hFFFF;
            12'd1023: out = 16'hFFFF;
            12'd1024: out = 16'hFFFF;
            12'd1025: out = 16'hFFC0;
            12'd1026: out = 16'hFF80;
            12'd1027: out = 16'hFF41;
            12'd1028: out = 16'hFF01;
            12'd1029: out = 16'hFEC2;
            12'd1030: out = 16'hFE82;
            12'd1031: out = 16'hFE43;
            12'd1032: out = 16'hFE04;
            12'd1033: out = 16'hFDC5;
            12'd1034: out = 16'hFD86;
            12'd1035: out = 16'hFD47;
            12'd1036: out = 16'hFD09;
            12'd1037: out = 16'hFCCA;
            12'd1038: out = 16'hFC8C;
            12'd1039: out = 16'hFC4E;
            12'd1040: out = 16'hFC10;
            12'd1041: out = 16'hFBD2;
            12'd1042: out = 16'hFB94;
            12'd1043: out = 16'hFB56;
            12'd1044: out = 16'hFB19;
            12'd1045: out = 16'hFADB;
            12'd1046: out = 16'hFA9E;
            12'd1047: out = 16'hFA60;
            12'd1048: out = 16'hFA23;
            12'd1049: out = 16'hF9E6;
            12'd1050: out = 16'hF9A9;
            12'd1051: out = 16'hF96C;
            12'd1052: out = 16'hF930;
            12'd1053: out = 16'hF8F3;
            12'd1054: out = 16'hF8B7;
            12'd1055: out = 16'hF87A;
            12'd1056: out = 16'hF83E;
            12'd1057: out = 16'hF802;
            12'd1058: out = 16'hF7C6;
            12'd1059: out = 16'hF78A;
            12'd1060: out = 16'hF74E;
            12'd1061: out = 16'hF713;
            12'd1062: out = 16'hF6D7;
            12'd1063: out = 16'hF69C;
            12'd1064: out = 16'hF660;
            12'd1065: out = 16'hF625;
            12'd1066: out = 16'hF5EA;
            12'd1067: out = 16'hF5AF;
            12'd1068: out = 16'hF574;
            12'd1069: out = 16'hF539;
            12'd1070: out = 16'hF4FF;
            12'd1071: out = 16'hF4C4;
            12'd1072: out = 16'hF48A;
            12'd1073: out = 16'hF44F;
            12'd1074: out = 16'hF415;
            12'd1075: out = 16'hF3DB;
            12'd1076: out = 16'hF3A1;
            12'd1077: out = 16'hF367;
            12'd1078: out = 16'hF32D;
            12'd1079: out = 16'hF2F3;
            12'd1080: out = 16'hF2BA;
            12'd1081: out = 16'hF280;
            12'd1082: out = 16'hF247;
            12'd1083: out = 16'hF20E;
            12'd1084: out = 16'hF1D5;
            12'd1085: out = 16'hF19B;
            12'd1086: out = 16'hF163;
            12'd1087: out = 16'hF12A;
            12'd1088: out = 16'hF0F1;
            12'd1089: out = 16'hF0B8;
            12'd1090: out = 16'hF080;
            12'd1091: out = 16'hF047;
            12'd1092: out = 16'hF00F;
            12'd1093: out = 16'hEFD7;
            12'd1094: out = 16'hEF9F;
            12'd1095: out = 16'hEF67;
            12'd1096: out = 16'hEF2F;
            12'd1097: out = 16'hEEF7;
            12'd1098: out = 16'hEEBF;
            12'd1099: out = 16'hEE88;
            12'd1100: out = 16'hEE50;
            12'd1101: out = 16'hEE19;
            12'd1102: out = 16'hEDE1;
            12'd1103: out = 16'hEDAA;
            12'd1104: out = 16'hED73;
            12'd1105: out = 16'hED3C;
            12'd1106: out = 16'hED05;
            12'd1107: out = 16'hECCE;
            12'd1108: out = 16'hEC98;
            12'd1109: out = 16'hEC61;
            12'd1110: out = 16'hEC2A;
            12'd1111: out = 16'hEBF4;
            12'd1112: out = 16'hEBBE;
            12'd1113: out = 16'hEB87;
            12'd1114: out = 16'hEB51;
            12'd1115: out = 16'hEB1B;
            12'd1116: out = 16'hEAE5;
            12'd1117: out = 16'hEAB0;
            12'd1118: out = 16'hEA7A;
            12'd1119: out = 16'hEA44;
            12'd1120: out = 16'hEA0F;
            12'd1121: out = 16'hE9D9;
            12'd1122: out = 16'hE9A4;
            12'd1123: out = 16'hE96F;
            12'd1124: out = 16'hE939;
            12'd1125: out = 16'hE904;
            12'd1126: out = 16'hE8CF;
            12'd1127: out = 16'hE89A;
            12'd1128: out = 16'hE866;
            12'd1129: out = 16'hE831;
            12'd1130: out = 16'hE7FC;
            12'd1131: out = 16'hE7C8;
            12'd1132: out = 16'hE793;
            12'd1133: out = 16'hE75F;
            12'd1134: out = 16'hE72B;
            12'd1135: out = 16'hE6F7;
            12'd1136: out = 16'hE6C3;
            12'd1137: out = 16'hE68F;
            12'd1138: out = 16'hE65B;
            12'd1139: out = 16'hE627;
            12'd1140: out = 16'hE5F3;
            12'd1141: out = 16'hE5C0;
            12'd1142: out = 16'hE58C;
            12'd1143: out = 16'hE559;
            12'd1144: out = 16'hE526;
            12'd1145: out = 16'hE4F2;
            12'd1146: out = 16'hE4BF;
            12'd1147: out = 16'hE48C;
            12'd1148: out = 16'hE459;
            12'd1149: out = 16'hE426;
            12'd1150: out = 16'hE3F4;
            12'd1151: out = 16'hE3C1;
            12'd1152: out = 16'hE38E;
            12'd1153: out = 16'hE35C;
            12'd1154: out = 16'hE329;
            12'd1155: out = 16'hE2F7;
            12'd1156: out = 16'hE2C5;
            12'd1157: out = 16'hE292;
            12'd1158: out = 16'hE260;
            12'd1159: out = 16'hE22E;
            12'd1160: out = 16'hE1FC;
            12'd1161: out = 16'hE1CB;
            12'd1162: out = 16'hE199;
            12'd1163: out = 16'hE167;
            12'd1164: out = 16'hE136;
            12'd1165: out = 16'hE104;
            12'd1166: out = 16'hE0D3;
            12'd1167: out = 16'hE0A1;
            12'd1168: out = 16'hE070;
            12'd1169: out = 16'hE03F;
            12'd1170: out = 16'hE00E;
            12'd1171: out = 16'hDFDD;
            12'd1172: out = 16'hDFAC;
            12'd1173: out = 16'hDF7B;
            12'd1174: out = 16'hDF4B;
            12'd1175: out = 16'hDF1A;
            12'd1176: out = 16'hDEE9;
            12'd1177: out = 16'hDEB9;
            12'd1178: out = 16'hDE88;
            12'd1179: out = 16'hDE58;
            12'd1180: out = 16'hDE28;
            12'd1181: out = 16'hDDF8;
            12'd1182: out = 16'hDDC8;
            12'd1183: out = 16'hDD98;
            12'd1184: out = 16'hDD68;
            12'd1185: out = 16'hDD38;
            12'd1186: out = 16'hDD08;
            12'd1187: out = 16'hDCD9;
            12'd1188: out = 16'hDCA9;
            12'd1189: out = 16'hDC79;
            12'd1190: out = 16'hDC4A;
            12'd1191: out = 16'hDC1B;
            12'd1192: out = 16'hDBEB;
            12'd1193: out = 16'hDBBC;
            12'd1194: out = 16'hDB8D;
            12'd1195: out = 16'hDB5E;
            12'd1196: out = 16'hDB2F;
            12'd1197: out = 16'hDB00;
            12'd1198: out = 16'hDAD1;
            12'd1199: out = 16'hDAA3;
            12'd1200: out = 16'hDA74;
            12'd1201: out = 16'hDA45;
            12'd1202: out = 16'hDA17;
            12'd1203: out = 16'hD9E9;
            12'd1204: out = 16'hD9BA;
            12'd1205: out = 16'hD98C;
            12'd1206: out = 16'hD95E;
            12'd1207: out = 16'hD930;
            12'd1208: out = 16'hD902;
            12'd1209: out = 16'hD8D4;
            12'd1210: out = 16'hD8A6;
            12'd1211: out = 16'hD878;
            12'd1212: out = 16'hD84A;
            12'd1213: out = 16'hD81D;
            12'd1214: out = 16'hD7EF;
            12'd1215: out = 16'hD7C2;
            12'd1216: out = 16'hD794;
            12'd1217: out = 16'hD767;
            12'd1218: out = 16'hD73A;
            12'd1219: out = 16'hD70C;
            12'd1220: out = 16'hD6DF;
            12'd1221: out = 16'hD6B2;
            12'd1222: out = 16'hD685;
            12'd1223: out = 16'hD658;
            12'd1224: out = 16'hD62C;
            12'd1225: out = 16'hD5FF;
            12'd1226: out = 16'hD5D2;
            12'd1227: out = 16'hD5A5;
            12'd1228: out = 16'hD579;
            12'd1229: out = 16'hD54C;
            12'd1230: out = 16'hD520;
            12'd1231: out = 16'hD4F4;
            12'd1232: out = 16'hD4C7;
            12'd1233: out = 16'hD49B;
            12'd1234: out = 16'hD46F;
            12'd1235: out = 16'hD443;
            12'd1236: out = 16'hD417;
            12'd1237: out = 16'hD3EB;
            12'd1238: out = 16'hD3BF;
            12'd1239: out = 16'hD394;
            12'd1240: out = 16'hD368;
            12'd1241: out = 16'hD33C;
            12'd1242: out = 16'hD311;
            12'd1243: out = 16'hD2E5;
            12'd1244: out = 16'hD2BA;
            12'd1245: out = 16'hD28F;
            12'd1246: out = 16'hD263;
            12'd1247: out = 16'hD238;
            12'd1248: out = 16'hD20D;
            12'd1249: out = 16'hD1E2;
            12'd1250: out = 16'hD1B7;
            12'd1251: out = 16'hD18C;
            12'd1252: out = 16'hD161;
            12'd1253: out = 16'hD137;
            12'd1254: out = 16'hD10C;
            12'd1255: out = 16'hD0E1;
            12'd1256: out = 16'hD0B7;
            12'd1257: out = 16'hD08C;
            12'd1258: out = 16'hD062;
            12'd1259: out = 16'hD037;
            12'd1260: out = 16'hD00D;
            12'd1261: out = 16'hCFE3;
            12'd1262: out = 16'hCFB9;
            12'd1263: out = 16'hCF8E;
            12'd1264: out = 16'hCF64;
            12'd1265: out = 16'hCF3A;
            12'd1266: out = 16'hCF11;
            12'd1267: out = 16'hCEE7;
            12'd1268: out = 16'hCEBD;
            12'd1269: out = 16'hCE93;
            12'd1270: out = 16'hCE6A;
            12'd1271: out = 16'hCE40;
            12'd1272: out = 16'hCE17;
            12'd1273: out = 16'hCDED;
            12'd1274: out = 16'hCDC4;
            12'd1275: out = 16'hCD9A;
            12'd1276: out = 16'hCD71;
            12'd1277: out = 16'hCD48;
            12'd1278: out = 16'hCD1F;
            12'd1279: out = 16'hCCF6;
            12'd1280: out = 16'hCCCD;
            12'd1281: out = 16'hCCA4;
            12'd1282: out = 16'hCC7B;
            12'd1283: out = 16'hCC52;
            12'd1284: out = 16'hCC29;
            12'd1285: out = 16'hCC01;
            12'd1286: out = 16'hCBD8;
            12'd1287: out = 16'hCBB0;
            12'd1288: out = 16'hCB87;
            12'd1289: out = 16'hCB5F;
            12'd1290: out = 16'hCB36;
            12'd1291: out = 16'hCB0E;
            12'd1292: out = 16'hCAE6;
            12'd1293: out = 16'hCABE;
            12'd1294: out = 16'hCA96;
            12'd1295: out = 16'hCA6E;
            12'd1296: out = 16'hCA46;
            12'd1297: out = 16'hCA1E;
            12'd1298: out = 16'hC9F6;
            12'd1299: out = 16'hC9CE;
            12'd1300: out = 16'hC9A6;
            12'd1301: out = 16'hC97F;
            12'd1302: out = 16'hC957;
            12'd1303: out = 16'hC92F;
            12'd1304: out = 16'hC908;
            12'd1305: out = 16'hC8E0;
            12'd1306: out = 16'hC8B9;
            12'd1307: out = 16'hC892;
            12'd1308: out = 16'hC86A;
            12'd1309: out = 16'hC843;
            12'd1310: out = 16'hC81C;
            12'd1311: out = 16'hC7F5;
            12'd1312: out = 16'hC7CE;
            12'd1313: out = 16'hC7A7;
            12'd1314: out = 16'hC780;
            12'd1315: out = 16'hC759;
            12'd1316: out = 16'hC733;
            12'd1317: out = 16'hC70C;
            12'd1318: out = 16'hC6E5;
            12'd1319: out = 16'hC6BF;
            12'd1320: out = 16'hC698;
            12'd1321: out = 16'hC672;
            12'd1322: out = 16'hC64B;
            12'd1323: out = 16'hC625;
            12'd1324: out = 16'hC5FE;
            12'd1325: out = 16'hC5D8;
            12'd1326: out = 16'hC5B2;
            12'd1327: out = 16'hC58C;
            12'd1328: out = 16'hC566;
            12'd1329: out = 16'hC540;
            12'd1330: out = 16'hC51A;
            12'd1331: out = 16'hC4F4;
            12'd1332: out = 16'hC4CE;
            12'd1333: out = 16'hC4A8;
            12'd1334: out = 16'hC482;
            12'd1335: out = 16'hC45D;
            12'd1336: out = 16'hC437;
            12'd1337: out = 16'hC412;
            12'd1338: out = 16'hC3EC;
            12'd1339: out = 16'hC3C7;
            12'd1340: out = 16'hC3A1;
            12'd1341: out = 16'hC37C;
            12'd1342: out = 16'hC357;
            12'd1343: out = 16'hC331;
            12'd1344: out = 16'hC30C;
            12'd1345: out = 16'hC2E7;
            12'd1346: out = 16'hC2C2;
            12'd1347: out = 16'hC29D;
            12'd1348: out = 16'hC278;
            12'd1349: out = 16'hC253;
            12'd1350: out = 16'hC22E;
            12'd1351: out = 16'hC209;
            12'd1352: out = 16'hC1E5;
            12'd1353: out = 16'hC1C0;
            12'd1354: out = 16'hC19B;
            12'd1355: out = 16'hC177;
            12'd1356: out = 16'hC152;
            12'd1357: out = 16'hC12E;
            12'd1358: out = 16'hC109;
            12'd1359: out = 16'hC0E5;
            12'd1360: out = 16'hC0C1;
            12'd1361: out = 16'hC09C;
            12'd1362: out = 16'hC078;
            12'd1363: out = 16'hC054;
            12'd1364: out = 16'hC030;
            12'd1365: out = 16'hC00C;
            12'd1366: out = 16'hBFE8;
            12'd1367: out = 16'hBFC4;
            12'd1368: out = 16'hBFA0;
            12'd1369: out = 16'hBF7C;
            12'd1370: out = 16'hBF59;
            12'd1371: out = 16'hBF35;
            12'd1372: out = 16'hBF11;
            12'd1373: out = 16'hBEEE;
            12'd1374: out = 16'hBECA;
            12'd1375: out = 16'hBEA6;
            12'd1376: out = 16'hBE83;
            12'd1377: out = 16'hBE60;
            12'd1378: out = 16'hBE3C;
            12'd1379: out = 16'hBE19;
            12'd1380: out = 16'hBDF6;
            12'd1381: out = 16'hBDD2;
            12'd1382: out = 16'hBDAF;
            12'd1383: out = 16'hBD8C;
            12'd1384: out = 16'hBD69;
            12'd1385: out = 16'hBD46;
            12'd1386: out = 16'hBD23;
            12'd1387: out = 16'hBD00;
            12'd1388: out = 16'hBCDD;
            12'd1389: out = 16'hBCBB;
            12'd1390: out = 16'hBC98;
            12'd1391: out = 16'hBC75;
            12'd1392: out = 16'hBC52;
            12'd1393: out = 16'hBC30;
            12'd1394: out = 16'hBC0D;
            12'd1395: out = 16'hBBEB;
            12'd1396: out = 16'hBBC8;
            12'd1397: out = 16'hBBA6;
            12'd1398: out = 16'hBB83;
            12'd1399: out = 16'hBB61;
            12'd1400: out = 16'hBB3F;
            12'd1401: out = 16'hBB1D;
            12'd1402: out = 16'hBAFB;
            12'd1403: out = 16'hBAD8;
            12'd1404: out = 16'hBAB6;
            12'd1405: out = 16'hBA94;
            12'd1406: out = 16'hBA72;
            12'd1407: out = 16'hBA50;
            12'd1408: out = 16'hBA2F;
            12'd1409: out = 16'hBA0D;
            12'd1410: out = 16'hB9EB;
            12'd1411: out = 16'hB9C9;
            12'd1412: out = 16'hB9A8;
            12'd1413: out = 16'hB986;
            12'd1414: out = 16'hB964;
            12'd1415: out = 16'hB943;
            12'd1416: out = 16'hB921;
            12'd1417: out = 16'hB900;
            12'd1418: out = 16'hB8DE;
            12'd1419: out = 16'hB8BD;
            12'd1420: out = 16'hB89C;
            12'd1421: out = 16'hB87B;
            12'd1422: out = 16'hB859;
            12'd1423: out = 16'hB838;
            12'd1424: out = 16'hB817;
            12'd1425: out = 16'hB7F6;
            12'd1426: out = 16'hB7D5;
            12'd1427: out = 16'hB7B4;
            12'd1428: out = 16'hB793;
            12'd1429: out = 16'hB772;
            12'd1430: out = 16'hB751;
            12'd1431: out = 16'hB730;
            12'd1432: out = 16'hB710;
            12'd1433: out = 16'hB6EF;
            12'd1434: out = 16'hB6CE;
            12'd1435: out = 16'hB6AE;
            12'd1436: out = 16'hB68D;
            12'd1437: out = 16'hB66D;
            12'd1438: out = 16'hB64C;
            12'd1439: out = 16'hB62C;
            12'd1440: out = 16'hB60B;
            12'd1441: out = 16'hB5EB;
            12'd1442: out = 16'hB5CB;
            12'd1443: out = 16'hB5AA;
            12'd1444: out = 16'hB58A;
            12'd1445: out = 16'hB56A;
            12'd1446: out = 16'hB54A;
            12'd1447: out = 16'hB52A;
            12'd1448: out = 16'hB50A;
            12'd1449: out = 16'hB4EA;
            12'd1450: out = 16'hB4CA;
            12'd1451: out = 16'hB4AA;
            12'd1452: out = 16'hB48A;
            12'd1453: out = 16'hB46A;
            12'd1454: out = 16'hB44B;
            12'd1455: out = 16'hB42B;
            12'd1456: out = 16'hB40B;
            12'd1457: out = 16'hB3EC;
            12'd1458: out = 16'hB3CC;
            12'd1459: out = 16'hB3AC;
            12'd1460: out = 16'hB38D;
            12'd1461: out = 16'hB36E;
            12'd1462: out = 16'hB34E;
            12'd1463: out = 16'hB32F;
            12'd1464: out = 16'hB30F;
            12'd1465: out = 16'hB2F0;
            12'd1466: out = 16'hB2D1;
            12'd1467: out = 16'hB2B2;
            12'd1468: out = 16'hB292;
            12'd1469: out = 16'hB273;
            12'd1470: out = 16'hB254;
            12'd1471: out = 16'hB235;
            12'd1472: out = 16'hB216;
            12'd1473: out = 16'hB1F7;
            12'd1474: out = 16'hB1D8;
            12'd1475: out = 16'hB1BA;
            12'd1476: out = 16'hB19B;
            12'd1477: out = 16'hB17C;
            12'd1478: out = 16'hB15D;
            12'd1479: out = 16'hB13E;
            12'd1480: out = 16'hB120;
            12'd1481: out = 16'hB101;
            12'd1482: out = 16'hB0E3;
            12'd1483: out = 16'hB0C4;
            12'd1484: out = 16'hB0A6;
            12'd1485: out = 16'hB087;
            12'd1486: out = 16'hB069;
            12'd1487: out = 16'hB04A;
            12'd1488: out = 16'hB02C;
            12'd1489: out = 16'hB00E;
            12'd1490: out = 16'hAFF0;
            12'd1491: out = 16'hAFD1;
            12'd1492: out = 16'hAFB3;
            12'd1493: out = 16'hAF95;
            12'd1494: out = 16'hAF77;
            12'd1495: out = 16'hAF59;
            12'd1496: out = 16'hAF3B;
            12'd1497: out = 16'hAF1D;
            12'd1498: out = 16'hAEFF;
            12'd1499: out = 16'hAEE1;
            12'd1500: out = 16'hAEC3;
            12'd1501: out = 16'hAEA5;
            12'd1502: out = 16'hAE88;
            12'd1503: out = 16'hAE6A;
            12'd1504: out = 16'hAE4C;
            12'd1505: out = 16'hAE2F;
            12'd1506: out = 16'hAE11;
            12'd1507: out = 16'hADF3;
            12'd1508: out = 16'hADD6;
            12'd1509: out = 16'hADB8;
            12'd1510: out = 16'hAD9B;
            12'd1511: out = 16'hAD7E;
            12'd1512: out = 16'hAD60;
            12'd1513: out = 16'hAD43;
            12'd1514: out = 16'hAD26;
            12'd1515: out = 16'hAD08;
            12'd1516: out = 16'hACEB;
            12'd1517: out = 16'hACCE;
            12'd1518: out = 16'hACB1;
            12'd1519: out = 16'hAC94;
            12'd1520: out = 16'hAC77;
            12'd1521: out = 16'hAC5A;
            12'd1522: out = 16'hAC3D;
            12'd1523: out = 16'hAC20;
            12'd1524: out = 16'hAC03;
            12'd1525: out = 16'hABE6;
            12'd1526: out = 16'hABC9;
            12'd1527: out = 16'hABAC;
            12'd1528: out = 16'hAB8F;
            12'd1529: out = 16'hAB73;
            12'd1530: out = 16'hAB56;
            12'd1531: out = 16'hAB39;
            12'd1532: out = 16'hAB1D;
            12'd1533: out = 16'hAB00;
            12'd1534: out = 16'hAAE4;
            12'd1535: out = 16'hAAC7;
            12'd1536: out = 16'hAAAB;
            12'd1537: out = 16'hAA8E;
            12'd1538: out = 16'hAA72;
            12'd1539: out = 16'hAA55;
            12'd1540: out = 16'hAA39;
            12'd1541: out = 16'hAA1D;
            12'd1542: out = 16'hAA01;
            12'd1543: out = 16'hA9E4;
            12'd1544: out = 16'hA9C8;
            12'd1545: out = 16'hA9AC;
            12'd1546: out = 16'hA990;
            12'd1547: out = 16'hA974;
            12'd1548: out = 16'hA958;
            12'd1549: out = 16'hA93C;
            12'd1550: out = 16'hA920;
            12'd1551: out = 16'hA904;
            12'd1552: out = 16'hA8E8;
            12'd1553: out = 16'hA8CC;
            12'd1554: out = 16'hA8B1;
            12'd1555: out = 16'hA895;
            12'd1556: out = 16'hA879;
            12'd1557: out = 16'hA85D;
            12'd1558: out = 16'hA842;
            12'd1559: out = 16'hA826;
            12'd1560: out = 16'hA80B;
            12'd1561: out = 16'hA7EF;
            12'd1562: out = 16'hA7D3;
            12'd1563: out = 16'hA7B8;
            12'd1564: out = 16'hA79C;
            12'd1565: out = 16'hA781;
            12'd1566: out = 16'hA766;
            12'd1567: out = 16'hA74A;
            12'd1568: out = 16'hA72F;
            12'd1569: out = 16'hA714;
            12'd1570: out = 16'hA6F8;
            12'd1571: out = 16'hA6DD;
            12'd1572: out = 16'hA6C2;
            12'd1573: out = 16'hA6A7;
            12'd1574: out = 16'hA68C;
            12'd1575: out = 16'hA671;
            12'd1576: out = 16'hA656;
            12'd1577: out = 16'hA63B;
            12'd1578: out = 16'hA620;
            12'd1579: out = 16'hA605;
            12'd1580: out = 16'hA5EA;
            12'd1581: out = 16'hA5CF;
            12'd1582: out = 16'hA5B4;
            12'd1583: out = 16'hA599;
            12'd1584: out = 16'hA57F;
            12'd1585: out = 16'hA564;
            12'd1586: out = 16'hA549;
            12'd1587: out = 16'hA52F;
            12'd1588: out = 16'hA514;
            12'd1589: out = 16'hA4F9;
            12'd1590: out = 16'hA4DF;
            12'd1591: out = 16'hA4C4;
            12'd1592: out = 16'hA4AA;
            12'd1593: out = 16'hA48F;
            12'd1594: out = 16'hA475;
            12'd1595: out = 16'hA45B;
            12'd1596: out = 16'hA440;
            12'd1597: out = 16'hA426;
            12'd1598: out = 16'hA40C;
            12'd1599: out = 16'hA3F1;
            12'd1600: out = 16'hA3D7;
            12'd1601: out = 16'hA3BD;
            12'd1602: out = 16'hA3A3;
            12'd1603: out = 16'hA389;
            12'd1604: out = 16'hA36E;
            12'd1605: out = 16'hA354;
            12'd1606: out = 16'hA33A;
            12'd1607: out = 16'hA320;
            12'd1608: out = 16'hA306;
            12'd1609: out = 16'hA2EC;
            12'd1610: out = 16'hA2D3;
            12'd1611: out = 16'hA2B9;
            12'd1612: out = 16'hA29F;
            12'd1613: out = 16'hA285;
            12'd1614: out = 16'hA26B;
            12'd1615: out = 16'hA251;
            12'd1616: out = 16'hA238;
            12'd1617: out = 16'hA21E;
            12'd1618: out = 16'hA204;
            12'd1619: out = 16'hA1EB;
            12'd1620: out = 16'hA1D1;
            12'd1621: out = 16'hA1B8;
            12'd1622: out = 16'hA19E;
            12'd1623: out = 16'hA185;
            12'd1624: out = 16'hA16B;
            12'd1625: out = 16'hA152;
            12'd1626: out = 16'hA138;
            12'd1627: out = 16'hA11F;
            12'd1628: out = 16'hA106;
            12'd1629: out = 16'hA0EC;
            12'd1630: out = 16'hA0D3;
            12'd1631: out = 16'hA0BA;
            12'd1632: out = 16'hA0A1;
            12'd1633: out = 16'hA087;
            12'd1634: out = 16'hA06E;
            12'd1635: out = 16'hA055;
            12'd1636: out = 16'hA03C;
            12'd1637: out = 16'hA023;
            12'd1638: out = 16'hA00A;
            12'd1639: out = 16'h9FF1;
            12'd1640: out = 16'h9FD8;
            12'd1641: out = 16'h9FBF;
            12'd1642: out = 16'h9FA6;
            12'd1643: out = 16'h9F8D;
            12'd1644: out = 16'h9F74;
            12'd1645: out = 16'h9F5C;
            12'd1646: out = 16'h9F43;
            12'd1647: out = 16'h9F2A;
            12'd1648: out = 16'h9F11;
            12'd1649: out = 16'h9EF9;
            12'd1650: out = 16'h9EE0;
            12'd1651: out = 16'h9EC7;
            12'd1652: out = 16'h9EAF;
            12'd1653: out = 16'h9E96;
            12'd1654: out = 16'h9E7E;
            12'd1655: out = 16'h9E65;
            12'd1656: out = 16'h9E4D;
            12'd1657: out = 16'h9E34;
            12'd1658: out = 16'h9E1C;
            12'd1659: out = 16'h9E03;
            12'd1660: out = 16'h9DEB;
            12'd1661: out = 16'h9DD3;
            12'd1662: out = 16'h9DBA;
            12'd1663: out = 16'h9DA2;
            12'd1664: out = 16'h9D8A;
            12'd1665: out = 16'h9D72;
            12'd1666: out = 16'h9D59;
            12'd1667: out = 16'h9D41;
            12'd1668: out = 16'h9D29;
            12'd1669: out = 16'h9D11;
            12'd1670: out = 16'h9CF9;
            12'd1671: out = 16'h9CE1;
            12'd1672: out = 16'h9CC9;
            12'd1673: out = 16'h9CB1;
            12'd1674: out = 16'h9C99;
            12'd1675: out = 16'h9C81;
            12'd1676: out = 16'h9C69;
            12'd1677: out = 16'h9C51;
            12'd1678: out = 16'h9C39;
            12'd1679: out = 16'h9C22;
            12'd1680: out = 16'h9C0A;
            12'd1681: out = 16'h9BF2;
            12'd1682: out = 16'h9BDA;
            12'd1683: out = 16'h9BC3;
            12'd1684: out = 16'h9BAB;
            12'd1685: out = 16'h9B93;
            12'd1686: out = 16'h9B7C;
            12'd1687: out = 16'h9B64;
            12'd1688: out = 16'h9B4C;
            12'd1689: out = 16'h9B35;
            12'd1690: out = 16'h9B1D;
            12'd1691: out = 16'h9B06;
            12'd1692: out = 16'h9AEE;
            12'd1693: out = 16'h9AD7;
            12'd1694: out = 16'h9AC0;
            12'd1695: out = 16'h9AA8;
            12'd1696: out = 16'h9A91;
            12'd1697: out = 16'h9A7A;
            12'd1698: out = 16'h9A62;
            12'd1699: out = 16'h9A4B;
            12'd1700: out = 16'h9A34;
            12'd1701: out = 16'h9A1D;
            12'd1702: out = 16'h9A05;
            12'd1703: out = 16'h99EE;
            12'd1704: out = 16'h99D7;
            12'd1705: out = 16'h99C0;
            12'd1706: out = 16'h99A9;
            12'd1707: out = 16'h9992;
            12'd1708: out = 16'h997B;
            12'd1709: out = 16'h9964;
            12'd1710: out = 16'h994D;
            12'd1711: out = 16'h9936;
            12'd1712: out = 16'h991F;
            12'd1713: out = 16'h9908;
            12'd1714: out = 16'h98F1;
            12'd1715: out = 16'h98DB;
            12'd1716: out = 16'h98C4;
            12'd1717: out = 16'h98AD;
            12'd1718: out = 16'h9896;
            12'd1719: out = 16'h987F;
            12'd1720: out = 16'h9869;
            12'd1721: out = 16'h9852;
            12'd1722: out = 16'h983B;
            12'd1723: out = 16'h9825;
            12'd1724: out = 16'h980E;
            12'd1725: out = 16'h97F8;
            12'd1726: out = 16'h97E1;
            12'd1727: out = 16'h97CB;
            12'd1728: out = 16'h97B4;
            12'd1729: out = 16'h979E;
            12'd1730: out = 16'h9787;
            12'd1731: out = 16'h9771;
            12'd1732: out = 16'h975A;
            12'd1733: out = 16'h9744;
            12'd1734: out = 16'h972E;
            12'd1735: out = 16'h9717;
            12'd1736: out = 16'h9701;
            12'd1737: out = 16'h96EB;
            12'd1738: out = 16'h96D5;
            12'd1739: out = 16'h96BE;
            12'd1740: out = 16'h96A8;
            12'd1741: out = 16'h9692;
            12'd1742: out = 16'h967C;
            12'd1743: out = 16'h9666;
            12'd1744: out = 16'h9650;
            12'd1745: out = 16'h963A;
            12'd1746: out = 16'h9624;
            12'd1747: out = 16'h960E;
            12'd1748: out = 16'h95F8;
            12'd1749: out = 16'h95E2;
            12'd1750: out = 16'h95CC;
            12'd1751: out = 16'h95B6;
            12'd1752: out = 16'h95A0;
            12'd1753: out = 16'h958A;
            12'd1754: out = 16'h9574;
            12'd1755: out = 16'h955F;
            12'd1756: out = 16'h9549;
            12'd1757: out = 16'h9533;
            12'd1758: out = 16'h951D;
            12'd1759: out = 16'h9508;
            12'd1760: out = 16'h94F2;
            12'd1761: out = 16'h94DC;
            12'd1762: out = 16'h94C7;
            12'd1763: out = 16'h94B1;
            12'd1764: out = 16'h949C;
            12'd1765: out = 16'h9486;
            12'd1766: out = 16'h9470;
            12'd1767: out = 16'h945B;
            12'd1768: out = 16'h9446;
            12'd1769: out = 16'h9430;
            12'd1770: out = 16'h941B;
            12'd1771: out = 16'h9405;
            12'd1772: out = 16'h93F0;
            12'd1773: out = 16'h93DA;
            12'd1774: out = 16'h93C5;
            12'd1775: out = 16'h93B0;
            12'd1776: out = 16'h939B;
            12'd1777: out = 16'h9385;
            12'd1778: out = 16'h9370;
            12'd1779: out = 16'h935B;
            12'd1780: out = 16'h9346;
            12'd1781: out = 16'h9330;
            12'd1782: out = 16'h931B;
            12'd1783: out = 16'h9306;
            12'd1784: out = 16'h92F1;
            12'd1785: out = 16'h92DC;
            12'd1786: out = 16'h92C7;
            12'd1787: out = 16'h92B2;
            12'd1788: out = 16'h929D;
            12'd1789: out = 16'h9288;
            12'd1790: out = 16'h9273;
            12'd1791: out = 16'h925E;
            12'd1792: out = 16'h9249;
            12'd1793: out = 16'h9234;
            12'd1794: out = 16'h921F;
            12'd1795: out = 16'h920B;
            12'd1796: out = 16'h91F6;
            12'd1797: out = 16'h91E1;
            12'd1798: out = 16'h91CC;
            12'd1799: out = 16'h91B7;
            12'd1800: out = 16'h91A3;
            12'd1801: out = 16'h918E;
            12'd1802: out = 16'h9179;
            12'd1803: out = 16'h9165;
            12'd1804: out = 16'h9150;
            12'd1805: out = 16'h913B;
            12'd1806: out = 16'h9127;
            12'd1807: out = 16'h9112;
            12'd1808: out = 16'h90FE;
            12'd1809: out = 16'h90E9;
            12'd1810: out = 16'h90D5;
            12'd1811: out = 16'h90C0;
            12'd1812: out = 16'h90AC;
            12'd1813: out = 16'h9097;
            12'd1814: out = 16'h9083;
            12'd1815: out = 16'h906F;
            12'd1816: out = 16'h905A;
            12'd1817: out = 16'h9046;
            12'd1818: out = 16'h9032;
            12'd1819: out = 16'h901D;
            12'd1820: out = 16'h9009;
            12'd1821: out = 16'h8FF5;
            12'd1822: out = 16'h8FE1;
            12'd1823: out = 16'h8FCC;
            12'd1824: out = 16'h8FB8;
            12'd1825: out = 16'h8FA4;
            12'd1826: out = 16'h8F90;
            12'd1827: out = 16'h8F7C;
            12'd1828: out = 16'h8F68;
            12'd1829: out = 16'h8F54;
            12'd1830: out = 16'h8F40;
            12'd1831: out = 16'h8F2B;
            12'd1832: out = 16'h8F17;
            12'd1833: out = 16'h8F03;
            12'd1834: out = 16'h8EF0;
            12'd1835: out = 16'h8EDC;
            12'd1836: out = 16'h8EC8;
            12'd1837: out = 16'h8EB4;
            12'd1838: out = 16'h8EA0;
            12'd1839: out = 16'h8E8C;
            12'd1840: out = 16'h8E78;
            12'd1841: out = 16'h8E64;
            12'd1842: out = 16'h8E51;
            12'd1843: out = 16'h8E3D;
            12'd1844: out = 16'h8E29;
            12'd1845: out = 16'h8E15;
            12'd1846: out = 16'h8E02;
            12'd1847: out = 16'h8DEE;
            12'd1848: out = 16'h8DDA;
            12'd1849: out = 16'h8DC7;
            12'd1850: out = 16'h8DB3;
            12'd1851: out = 16'h8D9F;
            12'd1852: out = 16'h8D8C;
            12'd1853: out = 16'h8D78;
            12'd1854: out = 16'h8D65;
            12'd1855: out = 16'h8D51;
            12'd1856: out = 16'h8D3E;
            12'd1857: out = 16'h8D2A;
            12'd1858: out = 16'h8D17;
            12'd1859: out = 16'h8D03;
            12'd1860: out = 16'h8CF0;
            12'd1861: out = 16'h8CDD;
            12'd1862: out = 16'h8CC9;
            12'd1863: out = 16'h8CB6;
            12'd1864: out = 16'h8CA3;
            12'd1865: out = 16'h8C8F;
            12'd1866: out = 16'h8C7C;
            12'd1867: out = 16'h8C69;
            12'd1868: out = 16'h8C56;
            12'd1869: out = 16'h8C42;
            12'd1870: out = 16'h8C2F;
            12'd1871: out = 16'h8C1C;
            12'd1872: out = 16'h8C09;
            12'd1873: out = 16'h8BF6;
            12'd1874: out = 16'h8BE2;
            12'd1875: out = 16'h8BCF;
            12'd1876: out = 16'h8BBC;
            12'd1877: out = 16'h8BA9;
            12'd1878: out = 16'h8B96;
            12'd1879: out = 16'h8B83;
            12'd1880: out = 16'h8B70;
            12'd1881: out = 16'h8B5D;
            12'd1882: out = 16'h8B4A;
            12'd1883: out = 16'h8B37;
            12'd1884: out = 16'h8B24;
            12'd1885: out = 16'h8B12;
            12'd1886: out = 16'h8AFF;
            12'd1887: out = 16'h8AEC;
            12'd1888: out = 16'h8AD9;
            12'd1889: out = 16'h8AC6;
            12'd1890: out = 16'h8AB3;
            12'd1891: out = 16'h8AA1;
            12'd1892: out = 16'h8A8E;
            12'd1893: out = 16'h8A7B;
            12'd1894: out = 16'h8A68;
            12'd1895: out = 16'h8A56;
            12'd1896: out = 16'h8A43;
            12'd1897: out = 16'h8A30;
            12'd1898: out = 16'h8A1E;
            12'd1899: out = 16'h8A0B;
            12'd1900: out = 16'h89F8;
            12'd1901: out = 16'h89E6;
            12'd1902: out = 16'h89D3;
            12'd1903: out = 16'h89C1;
            12'd1904: out = 16'h89AE;
            12'd1905: out = 16'h899C;
            12'd1906: out = 16'h8989;
            12'd1907: out = 16'h8977;
            12'd1908: out = 16'h8964;
            12'd1909: out = 16'h8952;
            12'd1910: out = 16'h8940;
            12'd1911: out = 16'h892D;
            12'd1912: out = 16'h891B;
            12'd1913: out = 16'h8908;
            12'd1914: out = 16'h88F6;
            12'd1915: out = 16'h88E4;
            12'd1916: out = 16'h88D2;
            12'd1917: out = 16'h88BF;
            12'd1918: out = 16'h88AD;
            12'd1919: out = 16'h889B;
            12'd1920: out = 16'h8889;
            12'd1921: out = 16'h8876;
            12'd1922: out = 16'h8864;
            12'd1923: out = 16'h8852;
            12'd1924: out = 16'h8840;
            12'd1925: out = 16'h882E;
            12'd1926: out = 16'h881C;
            12'd1927: out = 16'h880A;
            12'd1928: out = 16'h87F8;
            12'd1929: out = 16'h87E5;
            12'd1930: out = 16'h87D3;
            12'd1931: out = 16'h87C1;
            12'd1932: out = 16'h87AF;
            12'd1933: out = 16'h879D;
            12'd1934: out = 16'h878C;
            12'd1935: out = 16'h877A;
            12'd1936: out = 16'h8768;
            12'd1937: out = 16'h8756;
            12'd1938: out = 16'h8744;
            12'd1939: out = 16'h8732;
            12'd1940: out = 16'h8720;
            12'd1941: out = 16'h870E;
            12'd1942: out = 16'h86FD;
            12'd1943: out = 16'h86EB;
            12'd1944: out = 16'h86D9;
            12'd1945: out = 16'h86C7;
            12'd1946: out = 16'h86B6;
            12'd1947: out = 16'h86A4;
            12'd1948: out = 16'h8692;
            12'd1949: out = 16'h8680;
            12'd1950: out = 16'h866F;
            12'd1951: out = 16'h865D;
            12'd1952: out = 16'h864C;
            12'd1953: out = 16'h863A;
            12'd1954: out = 16'h8628;
            12'd1955: out = 16'h8617;
            12'd1956: out = 16'h8605;
            12'd1957: out = 16'h85F4;
            12'd1958: out = 16'h85E2;
            12'd1959: out = 16'h85D1;
            12'd1960: out = 16'h85BF;
            12'd1961: out = 16'h85AE;
            12'd1962: out = 16'h859C;
            12'd1963: out = 16'h858B;
            12'd1964: out = 16'h8579;
            12'd1965: out = 16'h8568;
            12'd1966: out = 16'h8557;
            12'd1967: out = 16'h8545;
            12'd1968: out = 16'h8534;
            12'd1969: out = 16'h8523;
            12'd1970: out = 16'h8511;
            12'd1971: out = 16'h8500;
            12'd1972: out = 16'h84EF;
            12'd1973: out = 16'h84DE;
            12'd1974: out = 16'h84CC;
            12'd1975: out = 16'h84BB;
            12'd1976: out = 16'h84AA;
            12'd1977: out = 16'h8499;
            12'd1978: out = 16'h8488;
            12'd1979: out = 16'h8476;
            12'd1980: out = 16'h8465;
            12'd1981: out = 16'h8454;
            12'd1982: out = 16'h8443;
            12'd1983: out = 16'h8432;
            12'd1984: out = 16'h8421;
            12'd1985: out = 16'h8410;
            12'd1986: out = 16'h83FF;
            12'd1987: out = 16'h83EE;
            12'd1988: out = 16'h83DD;
            12'd1989: out = 16'h83CC;
            12'd1990: out = 16'h83BB;
            12'd1991: out = 16'h83AA;
            12'd1992: out = 16'h8399;
            12'd1993: out = 16'h8388;
            12'd1994: out = 16'h8377;
            12'd1995: out = 16'h8367;
            12'd1996: out = 16'h8356;
            12'd1997: out = 16'h8345;
            12'd1998: out = 16'h8334;
            12'd1999: out = 16'h8323;
            12'd2000: out = 16'h8312;
            12'd2001: out = 16'h8302;
            12'd2002: out = 16'h82F1;
            12'd2003: out = 16'h82E0;
            12'd2004: out = 16'h82CF;
            12'd2005: out = 16'h82BF;
            12'd2006: out = 16'h82AE;
            12'd2007: out = 16'h829D;
            12'd2008: out = 16'h828D;
            12'd2009: out = 16'h827C;
            12'd2010: out = 16'h826B;
            12'd2011: out = 16'h825B;
            12'd2012: out = 16'h824A;
            12'd2013: out = 16'h823A;
            12'd2014: out = 16'h8229;
            12'd2015: out = 16'h8219;
            12'd2016: out = 16'h8208;
            12'd2017: out = 16'h81F8;
            12'd2018: out = 16'h81E7;
            12'd2019: out = 16'h81D7;
            12'd2020: out = 16'h81C6;
            12'd2021: out = 16'h81B6;
            12'd2022: out = 16'h81A5;
            12'd2023: out = 16'h8195;
            12'd2024: out = 16'h8185;
            12'd2025: out = 16'h8174;
            12'd2026: out = 16'h8164;
            12'd2027: out = 16'h8153;
            12'd2028: out = 16'h8143;
            12'd2029: out = 16'h8133;
            12'd2030: out = 16'h8123;
            12'd2031: out = 16'h8112;
            12'd2032: out = 16'h8102;
            12'd2033: out = 16'h80F2;
            12'd2034: out = 16'h80E2;
            12'd2035: out = 16'h80D1;
            12'd2036: out = 16'h80C1;
            12'd2037: out = 16'h80B1;
            12'd2038: out = 16'h80A1;
            12'd2039: out = 16'h8091;
            12'd2040: out = 16'h8081;
            12'd2041: out = 16'h8070;
            12'd2042: out = 16'h8060;
            12'd2043: out = 16'h8050;
            12'd2044: out = 16'h8040;
            12'd2045: out = 16'h8030;
            12'd2046: out = 16'h8020;
            12'd2047: out = 16'h8010;
            12'd2048: out = 16'h8000;
            12'd2049: out = 16'h7FF0;
            12'd2050: out = 16'h7FE0;
            12'd2051: out = 16'h7FD0;
            12'd2052: out = 16'h7FC0;
            12'd2053: out = 16'h7FB0;
            12'd2054: out = 16'h7FA0;
            12'd2055: out = 16'h7F90;
            12'd2056: out = 16'h7F80;
            12'd2057: out = 16'h7F71;
            12'd2058: out = 16'h7F61;
            12'd2059: out = 16'h7F51;
            12'd2060: out = 16'h7F41;
            12'd2061: out = 16'h7F31;
            12'd2062: out = 16'h7F22;
            12'd2063: out = 16'h7F12;
            12'd2064: out = 16'h7F02;
            12'd2065: out = 16'h7EF2;
            12'd2066: out = 16'h7EE3;
            12'd2067: out = 16'h7ED3;
            12'd2068: out = 16'h7EC3;
            12'd2069: out = 16'h7EB3;
            12'd2070: out = 16'h7EA4;
            12'd2071: out = 16'h7E94;
            12'd2072: out = 16'h7E84;
            12'd2073: out = 16'h7E75;
            12'd2074: out = 16'h7E65;
            12'd2075: out = 16'h7E56;
            12'd2076: out = 16'h7E46;
            12'd2077: out = 16'h7E36;
            12'd2078: out = 16'h7E27;
            12'd2079: out = 16'h7E17;
            12'd2080: out = 16'h7E08;
            12'd2081: out = 16'h7DF8;
            12'd2082: out = 16'h7DE9;
            12'd2083: out = 16'h7DD9;
            12'd2084: out = 16'h7DCA;
            12'd2085: out = 16'h7DBB;
            12'd2086: out = 16'h7DAB;
            12'd2087: out = 16'h7D9C;
            12'd2088: out = 16'h7D8C;
            12'd2089: out = 16'h7D7D;
            12'd2090: out = 16'h7D6E;
            12'd2091: out = 16'h7D5E;
            12'd2092: out = 16'h7D4F;
            12'd2093: out = 16'h7D3F;
            12'd2094: out = 16'h7D30;
            12'd2095: out = 16'h7D21;
            12'd2096: out = 16'h7D12;
            12'd2097: out = 16'h7D02;
            12'd2098: out = 16'h7CF3;
            12'd2099: out = 16'h7CE4;
            12'd2100: out = 16'h7CD5;
            12'd2101: out = 16'h7CC5;
            12'd2102: out = 16'h7CB6;
            12'd2103: out = 16'h7CA7;
            12'd2104: out = 16'h7C98;
            12'd2105: out = 16'h7C89;
            12'd2106: out = 16'h7C7A;
            12'd2107: out = 16'h7C6A;
            12'd2108: out = 16'h7C5B;
            12'd2109: out = 16'h7C4C;
            12'd2110: out = 16'h7C3D;
            12'd2111: out = 16'h7C2E;
            12'd2112: out = 16'h7C1F;
            12'd2113: out = 16'h7C10;
            12'd2114: out = 16'h7C01;
            12'd2115: out = 16'h7BF2;
            12'd2116: out = 16'h7BE3;
            12'd2117: out = 16'h7BD4;
            12'd2118: out = 16'h7BC5;
            12'd2119: out = 16'h7BB6;
            12'd2120: out = 16'h7BA7;
            12'd2121: out = 16'h7B98;
            12'd2122: out = 16'h7B89;
            12'd2123: out = 16'h7B7A;
            12'd2124: out = 16'h7B6C;
            12'd2125: out = 16'h7B5D;
            12'd2126: out = 16'h7B4E;
            12'd2127: out = 16'h7B3F;
            12'd2128: out = 16'h7B30;
            12'd2129: out = 16'h7B21;
            12'd2130: out = 16'h7B13;
            12'd2131: out = 16'h7B04;
            12'd2132: out = 16'h7AF5;
            12'd2133: out = 16'h7AE6;
            12'd2134: out = 16'h7AD7;
            12'd2135: out = 16'h7AC9;
            12'd2136: out = 16'h7ABA;
            12'd2137: out = 16'h7AAB;
            12'd2138: out = 16'h7A9D;
            12'd2139: out = 16'h7A8E;
            12'd2140: out = 16'h7A7F;
            12'd2141: out = 16'h7A71;
            12'd2142: out = 16'h7A62;
            12'd2143: out = 16'h7A53;
            12'd2144: out = 16'h7A45;
            12'd2145: out = 16'h7A36;
            12'd2146: out = 16'h7A28;
            12'd2147: out = 16'h7A19;
            12'd2148: out = 16'h7A0A;
            12'd2149: out = 16'h79FC;
            12'd2150: out = 16'h79ED;
            12'd2151: out = 16'h79DF;
            12'd2152: out = 16'h79D0;
            12'd2153: out = 16'h79C2;
            12'd2154: out = 16'h79B3;
            12'd2155: out = 16'h79A5;
            12'd2156: out = 16'h7997;
            12'd2157: out = 16'h7988;
            12'd2158: out = 16'h797A;
            12'd2159: out = 16'h796B;
            12'd2160: out = 16'h795D;
            12'd2161: out = 16'h794F;
            12'd2162: out = 16'h7940;
            12'd2163: out = 16'h7932;
            12'd2164: out = 16'h7923;
            12'd2165: out = 16'h7915;
            12'd2166: out = 16'h7907;
            12'd2167: out = 16'h78F9;
            12'd2168: out = 16'h78EA;
            12'd2169: out = 16'h78DC;
            12'd2170: out = 16'h78CE;
            12'd2171: out = 16'h78BF;
            12'd2172: out = 16'h78B1;
            12'd2173: out = 16'h78A3;
            12'd2174: out = 16'h7895;
            12'd2175: out = 16'h7887;
            12'd2176: out = 16'h7878;
            12'd2177: out = 16'h786A;
            12'd2178: out = 16'h785C;
            12'd2179: out = 16'h784E;
            12'd2180: out = 16'h7840;
            12'd2181: out = 16'h7832;
            12'd2182: out = 16'h7824;
            12'd2183: out = 16'h7816;
            12'd2184: out = 16'h7808;
            12'd2185: out = 16'h77F9;
            12'd2186: out = 16'h77EB;
            12'd2187: out = 16'h77DD;
            12'd2188: out = 16'h77CF;
            12'd2189: out = 16'h77C1;
            12'd2190: out = 16'h77B3;
            12'd2191: out = 16'h77A5;
            12'd2192: out = 16'h7797;
            12'd2193: out = 16'h7789;
            12'd2194: out = 16'h777B;
            12'd2195: out = 16'h776E;
            12'd2196: out = 16'h7760;
            12'd2197: out = 16'h7752;
            12'd2198: out = 16'h7744;
            12'd2199: out = 16'h7736;
            12'd2200: out = 16'h7728;
            12'd2201: out = 16'h771A;
            12'd2202: out = 16'h770C;
            12'd2203: out = 16'h76FE;
            12'd2204: out = 16'h76F1;
            12'd2205: out = 16'h76E3;
            12'd2206: out = 16'h76D5;
            12'd2207: out = 16'h76C7;
            12'd2208: out = 16'h76BA;
            12'd2209: out = 16'h76AC;
            12'd2210: out = 16'h769E;
            12'd2211: out = 16'h7690;
            12'd2212: out = 16'h7683;
            12'd2213: out = 16'h7675;
            12'd2214: out = 16'h7667;
            12'd2215: out = 16'h7659;
            12'd2216: out = 16'h764C;
            12'd2217: out = 16'h763E;
            12'd2218: out = 16'h7630;
            12'd2219: out = 16'h7623;
            12'd2220: out = 16'h7615;
            12'd2221: out = 16'h7608;
            12'd2222: out = 16'h75FA;
            12'd2223: out = 16'h75EC;
            12'd2224: out = 16'h75DF;
            12'd2225: out = 16'h75D1;
            12'd2226: out = 16'h75C4;
            12'd2227: out = 16'h75B6;
            12'd2228: out = 16'h75A9;
            12'd2229: out = 16'h759B;
            12'd2230: out = 16'h758E;
            12'd2231: out = 16'h7580;
            12'd2232: out = 16'h7573;
            12'd2233: out = 16'h7565;
            12'd2234: out = 16'h7558;
            12'd2235: out = 16'h754A;
            12'd2236: out = 16'h753D;
            12'd2237: out = 16'h752F;
            12'd2238: out = 16'h7522;
            12'd2239: out = 16'h7515;
            12'd2240: out = 16'h7507;
            12'd2241: out = 16'h74FA;
            12'd2242: out = 16'h74ED;
            12'd2243: out = 16'h74DF;
            12'd2244: out = 16'h74D2;
            12'd2245: out = 16'h74C5;
            12'd2246: out = 16'h74B7;
            12'd2247: out = 16'h74AA;
            12'd2248: out = 16'h749D;
            12'd2249: out = 16'h748F;
            12'd2250: out = 16'h7482;
            12'd2251: out = 16'h7475;
            12'd2252: out = 16'h7468;
            12'd2253: out = 16'h745A;
            12'd2254: out = 16'h744D;
            12'd2255: out = 16'h7440;
            12'd2256: out = 16'h7433;
            12'd2257: out = 16'h7426;
            12'd2258: out = 16'h7418;
            12'd2259: out = 16'h740B;
            12'd2260: out = 16'h73FE;
            12'd2261: out = 16'h73F1;
            12'd2262: out = 16'h73E4;
            12'd2263: out = 16'h73D7;
            12'd2264: out = 16'h73CA;
            12'd2265: out = 16'h73BD;
            12'd2266: out = 16'h73B0;
            12'd2267: out = 16'h73A2;
            12'd2268: out = 16'h7395;
            12'd2269: out = 16'h7388;
            12'd2270: out = 16'h737B;
            12'd2271: out = 16'h736E;
            12'd2272: out = 16'h7361;
            12'd2273: out = 16'h7354;
            12'd2274: out = 16'h7347;
            12'd2275: out = 16'h733A;
            12'd2276: out = 16'h732D;
            12'd2277: out = 16'h7320;
            12'd2278: out = 16'h7314;
            12'd2279: out = 16'h7307;
            12'd2280: out = 16'h72FA;
            12'd2281: out = 16'h72ED;
            12'd2282: out = 16'h72E0;
            12'd2283: out = 16'h72D3;
            12'd2284: out = 16'h72C6;
            12'd2285: out = 16'h72B9;
            12'd2286: out = 16'h72AC;
            12'd2287: out = 16'h72A0;
            12'd2288: out = 16'h7293;
            12'd2289: out = 16'h7286;
            12'd2290: out = 16'h7279;
            12'd2291: out = 16'h726C;
            12'd2292: out = 16'h7260;
            12'd2293: out = 16'h7253;
            12'd2294: out = 16'h7246;
            12'd2295: out = 16'h7239;
            12'd2296: out = 16'h722D;
            12'd2297: out = 16'h7220;
            12'd2298: out = 16'h7213;
            12'd2299: out = 16'h7206;
            12'd2300: out = 16'h71FA;
            12'd2301: out = 16'h71ED;
            12'd2302: out = 16'h71E0;
            12'd2303: out = 16'h71D4;
            12'd2304: out = 16'h71C7;
            12'd2305: out = 16'h71BA;
            12'd2306: out = 16'h71AE;
            12'd2307: out = 16'h71A1;
            12'd2308: out = 16'h7195;
            12'd2309: out = 16'h7188;
            12'd2310: out = 16'h717B;
            12'd2311: out = 16'h716F;
            12'd2312: out = 16'h7162;
            12'd2313: out = 16'h7156;
            12'd2314: out = 16'h7149;
            12'd2315: out = 16'h713D;
            12'd2316: out = 16'h7130;
            12'd2317: out = 16'h7124;
            12'd2318: out = 16'h7117;
            12'd2319: out = 16'h710B;
            12'd2320: out = 16'h70FE;
            12'd2321: out = 16'h70F2;
            12'd2322: out = 16'h70E5;
            12'd2323: out = 16'h70D9;
            12'd2324: out = 16'h70CC;
            12'd2325: out = 16'h70C0;
            12'd2326: out = 16'h70B4;
            12'd2327: out = 16'h70A7;
            12'd2328: out = 16'h709B;
            12'd2329: out = 16'h708E;
            12'd2330: out = 16'h7082;
            12'd2331: out = 16'h7076;
            12'd2332: out = 16'h7069;
            12'd2333: out = 16'h705D;
            12'd2334: out = 16'h7051;
            12'd2335: out = 16'h7044;
            12'd2336: out = 16'h7038;
            12'd2337: out = 16'h702C;
            12'd2338: out = 16'h7020;
            12'd2339: out = 16'h7013;
            12'd2340: out = 16'h7007;
            12'd2341: out = 16'h6FFB;
            12'd2342: out = 16'h6FEF;
            12'd2343: out = 16'h6FE2;
            12'd2344: out = 16'h6FD6;
            12'd2345: out = 16'h6FCA;
            12'd2346: out = 16'h6FBE;
            12'd2347: out = 16'h6FB1;
            12'd2348: out = 16'h6FA5;
            12'd2349: out = 16'h6F99;
            12'd2350: out = 16'h6F8D;
            12'd2351: out = 16'h6F81;
            12'd2352: out = 16'h6F75;
            12'd2353: out = 16'h6F69;
            12'd2354: out = 16'h6F5C;
            12'd2355: out = 16'h6F50;
            12'd2356: out = 16'h6F44;
            12'd2357: out = 16'h6F38;
            12'd2358: out = 16'h6F2C;
            12'd2359: out = 16'h6F20;
            12'd2360: out = 16'h6F14;
            12'd2361: out = 16'h6F08;
            12'd2362: out = 16'h6EFC;
            12'd2363: out = 16'h6EF0;
            12'd2364: out = 16'h6EE4;
            12'd2365: out = 16'h6ED8;
            12'd2366: out = 16'h6ECC;
            12'd2367: out = 16'h6EC0;
            12'd2368: out = 16'h6EB4;
            12'd2369: out = 16'h6EA8;
            12'd2370: out = 16'h6E9C;
            12'd2371: out = 16'h6E90;
            12'd2372: out = 16'h6E84;
            12'd2373: out = 16'h6E78;
            12'd2374: out = 16'h6E6C;
            12'd2375: out = 16'h6E60;
            12'd2376: out = 16'h6E54;
            12'd2377: out = 16'h6E49;
            12'd2378: out = 16'h6E3D;
            12'd2379: out = 16'h6E31;
            12'd2380: out = 16'h6E25;
            12'd2381: out = 16'h6E19;
            12'd2382: out = 16'h6E0D;
            12'd2383: out = 16'h6E02;
            12'd2384: out = 16'h6DF6;
            12'd2385: out = 16'h6DEA;
            12'd2386: out = 16'h6DDE;
            12'd2387: out = 16'h6DD2;
            12'd2388: out = 16'h6DC7;
            12'd2389: out = 16'h6DBB;
            12'd2390: out = 16'h6DAF;
            12'd2391: out = 16'h6DA3;
            12'd2392: out = 16'h6D98;
            12'd2393: out = 16'h6D8C;
            12'd2394: out = 16'h6D80;
            12'd2395: out = 16'h6D74;
            12'd2396: out = 16'h6D69;
            12'd2397: out = 16'h6D5D;
            12'd2398: out = 16'h6D51;
            12'd2399: out = 16'h6D46;
            12'd2400: out = 16'h6D3A;
            12'd2401: out = 16'h6D2E;
            12'd2402: out = 16'h6D23;
            12'd2403: out = 16'h6D17;
            12'd2404: out = 16'h6D0C;
            12'd2405: out = 16'h6D00;
            12'd2406: out = 16'h6CF4;
            12'd2407: out = 16'h6CE9;
            12'd2408: out = 16'h6CDD;
            12'd2409: out = 16'h6CD2;
            12'd2410: out = 16'h6CC6;
            12'd2411: out = 16'h6CBA;
            12'd2412: out = 16'h6CAF;
            12'd2413: out = 16'h6CA3;
            12'd2414: out = 16'h6C98;
            12'd2415: out = 16'h6C8C;
            12'd2416: out = 16'h6C81;
            12'd2417: out = 16'h6C75;
            12'd2418: out = 16'h6C6A;
            12'd2419: out = 16'h6C5E;
            12'd2420: out = 16'h6C53;
            12'd2421: out = 16'h6C47;
            12'd2422: out = 16'h6C3C;
            12'd2423: out = 16'h6C31;
            12'd2424: out = 16'h6C25;
            12'd2425: out = 16'h6C1A;
            12'd2426: out = 16'h6C0E;
            12'd2427: out = 16'h6C03;
            12'd2428: out = 16'h6BF8;
            12'd2429: out = 16'h6BEC;
            12'd2430: out = 16'h6BE1;
            12'd2431: out = 16'h6BD5;
            12'd2432: out = 16'h6BCA;
            12'd2433: out = 16'h6BBF;
            12'd2434: out = 16'h6BB3;
            12'd2435: out = 16'h6BA8;
            12'd2436: out = 16'h6B9D;
            12'd2437: out = 16'h6B91;
            12'd2438: out = 16'h6B86;
            12'd2439: out = 16'h6B7B;
            12'd2440: out = 16'h6B70;
            12'd2441: out = 16'h6B64;
            12'd2442: out = 16'h6B59;
            12'd2443: out = 16'h6B4E;
            12'd2444: out = 16'h6B43;
            12'd2445: out = 16'h6B37;
            12'd2446: out = 16'h6B2C;
            12'd2447: out = 16'h6B21;
            12'd2448: out = 16'h6B16;
            12'd2449: out = 16'h6B0B;
            12'd2450: out = 16'h6AFF;
            12'd2451: out = 16'h6AF4;
            12'd2452: out = 16'h6AE9;
            12'd2453: out = 16'h6ADE;
            12'd2454: out = 16'h6AD3;
            12'd2455: out = 16'h6AC8;
            12'd2456: out = 16'h6ABC;
            12'd2457: out = 16'h6AB1;
            12'd2458: out = 16'h6AA6;
            12'd2459: out = 16'h6A9B;
            12'd2460: out = 16'h6A90;
            12'd2461: out = 16'h6A85;
            12'd2462: out = 16'h6A7A;
            12'd2463: out = 16'h6A6F;
            12'd2464: out = 16'h6A64;
            12'd2465: out = 16'h6A59;
            12'd2466: out = 16'h6A4E;
            12'd2467: out = 16'h6A43;
            12'd2468: out = 16'h6A38;
            12'd2469: out = 16'h6A2D;
            12'd2470: out = 16'h6A22;
            12'd2471: out = 16'h6A17;
            12'd2472: out = 16'h6A0C;
            12'd2473: out = 16'h6A01;
            12'd2474: out = 16'h69F6;
            12'd2475: out = 16'h69EB;
            12'd2476: out = 16'h69E0;
            12'd2477: out = 16'h69D5;
            12'd2478: out = 16'h69CA;
            12'd2479: out = 16'h69BF;
            12'd2480: out = 16'h69B4;
            12'd2481: out = 16'h69A9;
            12'd2482: out = 16'h699E;
            12'd2483: out = 16'h6993;
            12'd2484: out = 16'h6988;
            12'd2485: out = 16'h697E;
            12'd2486: out = 16'h6973;
            12'd2487: out = 16'h6968;
            12'd2488: out = 16'h695D;
            12'd2489: out = 16'h6952;
            12'd2490: out = 16'h6947;
            12'd2491: out = 16'h693D;
            12'd2492: out = 16'h6932;
            12'd2493: out = 16'h6927;
            12'd2494: out = 16'h691C;
            12'd2495: out = 16'h6911;
            12'd2496: out = 16'h6907;
            12'd2497: out = 16'h68FC;
            12'd2498: out = 16'h68F1;
            12'd2499: out = 16'h68E6;
            12'd2500: out = 16'h68DC;
            12'd2501: out = 16'h68D1;
            12'd2502: out = 16'h68C6;
            12'd2503: out = 16'h68BB;
            12'd2504: out = 16'h68B1;
            12'd2505: out = 16'h68A6;
            12'd2506: out = 16'h689B;
            12'd2507: out = 16'h6891;
            12'd2508: out = 16'h6886;
            12'd2509: out = 16'h687B;
            12'd2510: out = 16'h6871;
            12'd2511: out = 16'h6866;
            12'd2512: out = 16'h685B;
            12'd2513: out = 16'h6851;
            12'd2514: out = 16'h6846;
            12'd2515: out = 16'h683B;
            12'd2516: out = 16'h6831;
            12'd2517: out = 16'h6826;
            12'd2518: out = 16'h681C;
            12'd2519: out = 16'h6811;
            12'd2520: out = 16'h6807;
            12'd2521: out = 16'h67FC;
            12'd2522: out = 16'h67F1;
            12'd2523: out = 16'h67E7;
            12'd2524: out = 16'h67DC;
            12'd2525: out = 16'h67D2;
            12'd2526: out = 16'h67C7;
            12'd2527: out = 16'h67BD;
            12'd2528: out = 16'h67B2;
            12'd2529: out = 16'h67A8;
            12'd2530: out = 16'h679D;
            12'd2531: out = 16'h6793;
            12'd2532: out = 16'h6788;
            12'd2533: out = 16'h677E;
            12'd2534: out = 16'h6773;
            12'd2535: out = 16'h6769;
            12'd2536: out = 16'h675E;
            12'd2537: out = 16'h6754;
            12'd2538: out = 16'h674A;
            12'd2539: out = 16'h673F;
            12'd2540: out = 16'h6735;
            12'd2541: out = 16'h672A;
            12'd2542: out = 16'h6720;
            12'd2543: out = 16'h6716;
            12'd2544: out = 16'h670B;
            12'd2545: out = 16'h6701;
            12'd2546: out = 16'h66F7;
            12'd2547: out = 16'h66EC;
            12'd2548: out = 16'h66E2;
            12'd2549: out = 16'h66D8;
            12'd2550: out = 16'h66CD;
            12'd2551: out = 16'h66C3;
            12'd2552: out = 16'h66B9;
            12'd2553: out = 16'h66AE;
            12'd2554: out = 16'h66A4;
            12'd2555: out = 16'h669A;
            12'd2556: out = 16'h668F;
            12'd2557: out = 16'h6685;
            12'd2558: out = 16'h667B;
            12'd2559: out = 16'h6671;
            12'd2560: out = 16'h6666;
            12'd2561: out = 16'h665C;
            12'd2562: out = 16'h6652;
            12'd2563: out = 16'h6648;
            12'd2564: out = 16'h663E;
            12'd2565: out = 16'h6633;
            12'd2566: out = 16'h6629;
            12'd2567: out = 16'h661F;
            12'd2568: out = 16'h6615;
            12'd2569: out = 16'h660B;
            12'd2570: out = 16'h6600;
            12'd2571: out = 16'h65F6;
            12'd2572: out = 16'h65EC;
            12'd2573: out = 16'h65E2;
            12'd2574: out = 16'h65D8;
            12'd2575: out = 16'h65CE;
            12'd2576: out = 16'h65C4;
            12'd2577: out = 16'h65B9;
            12'd2578: out = 16'h65AF;
            12'd2579: out = 16'h65A5;
            12'd2580: out = 16'h659B;
            12'd2581: out = 16'h6591;
            12'd2582: out = 16'h6587;
            12'd2583: out = 16'h657D;
            12'd2584: out = 16'h6573;
            12'd2585: out = 16'h6569;
            12'd2586: out = 16'h655F;
            12'd2587: out = 16'h6555;
            12'd2588: out = 16'h654B;
            12'd2589: out = 16'h6541;
            12'd2590: out = 16'h6537;
            12'd2591: out = 16'h652D;
            12'd2592: out = 16'h6523;
            12'd2593: out = 16'h6519;
            12'd2594: out = 16'h650F;
            12'd2595: out = 16'h6505;
            12'd2596: out = 16'h64FB;
            12'd2597: out = 16'h64F1;
            12'd2598: out = 16'h64E7;
            12'd2599: out = 16'h64DD;
            12'd2600: out = 16'h64D3;
            12'd2601: out = 16'h64C9;
            12'd2602: out = 16'h64BF;
            12'd2603: out = 16'h64B5;
            12'd2604: out = 16'h64AB;
            12'd2605: out = 16'h64A2;
            12'd2606: out = 16'h6498;
            12'd2607: out = 16'h648E;
            12'd2608: out = 16'h6484;
            12'd2609: out = 16'h647A;
            12'd2610: out = 16'h6470;
            12'd2611: out = 16'h6466;
            12'd2612: out = 16'h645D;
            12'd2613: out = 16'h6453;
            12'd2614: out = 16'h6449;
            12'd2615: out = 16'h643F;
            12'd2616: out = 16'h6435;
            12'd2617: out = 16'h642B;
            12'd2618: out = 16'h6422;
            12'd2619: out = 16'h6418;
            12'd2620: out = 16'h640E;
            12'd2621: out = 16'h6404;
            12'd2622: out = 16'h63FB;
            12'd2623: out = 16'h63F1;
            12'd2624: out = 16'h63E7;
            12'd2625: out = 16'h63DD;
            12'd2626: out = 16'h63D4;
            12'd2627: out = 16'h63CA;
            12'd2628: out = 16'h63C0;
            12'd2629: out = 16'h63B6;
            12'd2630: out = 16'h63AD;
            12'd2631: out = 16'h63A3;
            12'd2632: out = 16'h6399;
            12'd2633: out = 16'h6390;
            12'd2634: out = 16'h6386;
            12'd2635: out = 16'h637C;
            12'd2636: out = 16'h6373;
            12'd2637: out = 16'h6369;
            12'd2638: out = 16'h635F;
            12'd2639: out = 16'h6356;
            12'd2640: out = 16'h634C;
            12'd2641: out = 16'h6342;
            12'd2642: out = 16'h6339;
            12'd2643: out = 16'h632F;
            12'd2644: out = 16'h6326;
            12'd2645: out = 16'h631C;
            12'd2646: out = 16'h6312;
            12'd2647: out = 16'h6309;
            12'd2648: out = 16'h62FF;
            12'd2649: out = 16'h62F6;
            12'd2650: out = 16'h62EC;
            12'd2651: out = 16'h62E3;
            12'd2652: out = 16'h62D9;
            12'd2653: out = 16'h62CF;
            12'd2654: out = 16'h62C6;
            12'd2655: out = 16'h62BC;
            12'd2656: out = 16'h62B3;
            12'd2657: out = 16'h62A9;
            12'd2658: out = 16'h62A0;
            12'd2659: out = 16'h6296;
            12'd2660: out = 16'h628D;
            12'd2661: out = 16'h6283;
            12'd2662: out = 16'h627A;
            12'd2663: out = 16'h6270;
            12'd2664: out = 16'h6267;
            12'd2665: out = 16'h625E;
            12'd2666: out = 16'h6254;
            12'd2667: out = 16'h624B;
            12'd2668: out = 16'h6241;
            12'd2669: out = 16'h6238;
            12'd2670: out = 16'h622E;
            12'd2671: out = 16'h6225;
            12'd2672: out = 16'h621C;
            12'd2673: out = 16'h6212;
            12'd2674: out = 16'h6209;
            12'd2675: out = 16'h61FF;
            12'd2676: out = 16'h61F6;
            12'd2677: out = 16'h61ED;
            12'd2678: out = 16'h61E3;
            12'd2679: out = 16'h61DA;
            12'd2680: out = 16'h61D1;
            12'd2681: out = 16'h61C7;
            12'd2682: out = 16'h61BE;
            12'd2683: out = 16'h61B5;
            12'd2684: out = 16'h61AB;
            12'd2685: out = 16'h61A2;
            12'd2686: out = 16'h6199;
            12'd2687: out = 16'h618F;
            12'd2688: out = 16'h6186;
            12'd2689: out = 16'h617D;
            12'd2690: out = 16'h6174;
            12'd2691: out = 16'h616A;
            12'd2692: out = 16'h6161;
            12'd2693: out = 16'h6158;
            12'd2694: out = 16'h614E;
            12'd2695: out = 16'h6145;
            12'd2696: out = 16'h613C;
            12'd2697: out = 16'h6133;
            12'd2698: out = 16'h612A;
            12'd2699: out = 16'h6120;
            12'd2700: out = 16'h6117;
            12'd2701: out = 16'h610E;
            12'd2702: out = 16'h6105;
            12'd2703: out = 16'h60FC;
            12'd2704: out = 16'h60F2;
            12'd2705: out = 16'h60E9;
            12'd2706: out = 16'h60E0;
            12'd2707: out = 16'h60D7;
            12'd2708: out = 16'h60CE;
            12'd2709: out = 16'h60C5;
            12'd2710: out = 16'h60BB;
            12'd2711: out = 16'h60B2;
            12'd2712: out = 16'h60A9;
            12'd2713: out = 16'h60A0;
            12'd2714: out = 16'h6097;
            12'd2715: out = 16'h608E;
            12'd2716: out = 16'h6085;
            12'd2717: out = 16'h607C;
            12'd2718: out = 16'h6073;
            12'd2719: out = 16'h6069;
            12'd2720: out = 16'h6060;
            12'd2721: out = 16'h6057;
            12'd2722: out = 16'h604E;
            12'd2723: out = 16'h6045;
            12'd2724: out = 16'h603C;
            12'd2725: out = 16'h6033;
            12'd2726: out = 16'h602A;
            12'd2727: out = 16'h6021;
            12'd2728: out = 16'h6018;
            12'd2729: out = 16'h600F;
            12'd2730: out = 16'h6006;
            12'd2731: out = 16'h5FFD;
            12'd2732: out = 16'h5FF4;
            12'd2733: out = 16'h5FEB;
            12'd2734: out = 16'h5FE2;
            12'd2735: out = 16'h5FD9;
            12'd2736: out = 16'h5FD0;
            12'd2737: out = 16'h5FC7;
            12'd2738: out = 16'h5FBE;
            12'd2739: out = 16'h5FB5;
            12'd2740: out = 16'h5FAC;
            12'd2741: out = 16'h5FA3;
            12'd2742: out = 16'h5F9A;
            12'd2743: out = 16'h5F91;
            12'd2744: out = 16'h5F89;
            12'd2745: out = 16'h5F80;
            12'd2746: out = 16'h5F77;
            12'd2747: out = 16'h5F6E;
            12'd2748: out = 16'h5F65;
            12'd2749: out = 16'h5F5C;
            12'd2750: out = 16'h5F53;
            12'd2751: out = 16'h5F4A;
            12'd2752: out = 16'h5F41;
            12'd2753: out = 16'h5F39;
            12'd2754: out = 16'h5F30;
            12'd2755: out = 16'h5F27;
            12'd2756: out = 16'h5F1E;
            12'd2757: out = 16'h5F15;
            12'd2758: out = 16'h5F0C;
            12'd2759: out = 16'h5F04;
            12'd2760: out = 16'h5EFB;
            12'd2761: out = 16'h5EF2;
            12'd2762: out = 16'h5EE9;
            12'd2763: out = 16'h5EE0;
            12'd2764: out = 16'h5ED8;
            12'd2765: out = 16'h5ECF;
            12'd2766: out = 16'h5EC6;
            12'd2767: out = 16'h5EBD;
            12'd2768: out = 16'h5EB5;
            12'd2769: out = 16'h5EAC;
            12'd2770: out = 16'h5EA3;
            12'd2771: out = 16'h5E9A;
            12'd2772: out = 16'h5E92;
            12'd2773: out = 16'h5E89;
            12'd2774: out = 16'h5E80;
            12'd2775: out = 16'h5E77;
            12'd2776: out = 16'h5E6F;
            12'd2777: out = 16'h5E66;
            12'd2778: out = 16'h5E5D;
            12'd2779: out = 16'h5E55;
            12'd2780: out = 16'h5E4C;
            12'd2781: out = 16'h5E43;
            12'd2782: out = 16'h5E3B;
            12'd2783: out = 16'h5E32;
            12'd2784: out = 16'h5E29;
            12'd2785: out = 16'h5E21;
            12'd2786: out = 16'h5E18;
            12'd2787: out = 16'h5E0F;
            12'd2788: out = 16'h5E07;
            12'd2789: out = 16'h5DFE;
            12'd2790: out = 16'h5DF5;
            12'd2791: out = 16'h5DED;
            12'd2792: out = 16'h5DE4;
            12'd2793: out = 16'h5DDC;
            12'd2794: out = 16'h5DD3;
            12'd2795: out = 16'h5DCA;
            12'd2796: out = 16'h5DC2;
            12'd2797: out = 16'h5DB9;
            12'd2798: out = 16'h5DB1;
            12'd2799: out = 16'h5DA8;
            12'd2800: out = 16'h5D9F;
            12'd2801: out = 16'h5D97;
            12'd2802: out = 16'h5D8E;
            12'd2803: out = 16'h5D86;
            12'd2804: out = 16'h5D7D;
            12'd2805: out = 16'h5D75;
            12'd2806: out = 16'h5D6C;
            12'd2807: out = 16'h5D64;
            12'd2808: out = 16'h5D5B;
            12'd2809: out = 16'h5D53;
            12'd2810: out = 16'h5D4A;
            12'd2811: out = 16'h5D42;
            12'd2812: out = 16'h5D39;
            12'd2813: out = 16'h5D31;
            12'd2814: out = 16'h5D28;
            12'd2815: out = 16'h5D20;
            12'd2816: out = 16'h5D17;
            12'd2817: out = 16'h5D0F;
            12'd2818: out = 16'h5D06;
            12'd2819: out = 16'h5CFE;
            12'd2820: out = 16'h5CF5;
            12'd2821: out = 16'h5CED;
            12'd2822: out = 16'h5CE5;
            12'd2823: out = 16'h5CDC;
            12'd2824: out = 16'h5CD4;
            12'd2825: out = 16'h5CCB;
            12'd2826: out = 16'h5CC3;
            12'd2827: out = 16'h5CBB;
            12'd2828: out = 16'h5CB2;
            12'd2829: out = 16'h5CAA;
            12'd2830: out = 16'h5CA1;
            12'd2831: out = 16'h5C99;
            12'd2832: out = 16'h5C91;
            12'd2833: out = 16'h5C88;
            12'd2834: out = 16'h5C80;
            12'd2835: out = 16'h5C78;
            12'd2836: out = 16'h5C6F;
            12'd2837: out = 16'h5C67;
            12'd2838: out = 16'h5C5F;
            12'd2839: out = 16'h5C56;
            12'd2840: out = 16'h5C4E;
            12'd2841: out = 16'h5C46;
            12'd2842: out = 16'h5C3D;
            12'd2843: out = 16'h5C35;
            12'd2844: out = 16'h5C2D;
            12'd2845: out = 16'h5C24;
            12'd2846: out = 16'h5C1C;
            12'd2847: out = 16'h5C14;
            12'd2848: out = 16'h5C0C;
            12'd2849: out = 16'h5C03;
            12'd2850: out = 16'h5BFB;
            12'd2851: out = 16'h5BF3;
            12'd2852: out = 16'h5BEA;
            12'd2853: out = 16'h5BE2;
            12'd2854: out = 16'h5BDA;
            12'd2855: out = 16'h5BD2;
            12'd2856: out = 16'h5BCA;
            12'd2857: out = 16'h5BC1;
            12'd2858: out = 16'h5BB9;
            12'd2859: out = 16'h5BB1;
            12'd2860: out = 16'h5BA9;
            12'd2861: out = 16'h5BA0;
            12'd2862: out = 16'h5B98;
            12'd2863: out = 16'h5B90;
            12'd2864: out = 16'h5B88;
            12'd2865: out = 16'h5B80;
            12'd2866: out = 16'h5B78;
            12'd2867: out = 16'h5B6F;
            12'd2868: out = 16'h5B67;
            12'd2869: out = 16'h5B5F;
            12'd2870: out = 16'h5B57;
            12'd2871: out = 16'h5B4F;
            12'd2872: out = 16'h5B47;
            12'd2873: out = 16'h5B3E;
            12'd2874: out = 16'h5B36;
            12'd2875: out = 16'h5B2E;
            12'd2876: out = 16'h5B26;
            12'd2877: out = 16'h5B1E;
            12'd2878: out = 16'h5B16;
            12'd2879: out = 16'h5B0E;
            12'd2880: out = 16'h5B06;
            12'd2881: out = 16'h5AFE;
            12'd2882: out = 16'h5AF6;
            12'd2883: out = 16'h5AED;
            12'd2884: out = 16'h5AE5;
            12'd2885: out = 16'h5ADD;
            12'd2886: out = 16'h5AD5;
            12'd2887: out = 16'h5ACD;
            12'd2888: out = 16'h5AC5;
            12'd2889: out = 16'h5ABD;
            12'd2890: out = 16'h5AB5;
            12'd2891: out = 16'h5AAD;
            12'd2892: out = 16'h5AA5;
            12'd2893: out = 16'h5A9D;
            12'd2894: out = 16'h5A95;
            12'd2895: out = 16'h5A8D;
            12'd2896: out = 16'h5A85;
            12'd2897: out = 16'h5A7D;
            12'd2898: out = 16'h5A75;
            12'd2899: out = 16'h5A6D;
            12'd2900: out = 16'h5A65;
            12'd2901: out = 16'h5A5D;
            12'd2902: out = 16'h5A55;
            12'd2903: out = 16'h5A4D;
            12'd2904: out = 16'h5A45;
            12'd2905: out = 16'h5A3D;
            12'd2906: out = 16'h5A35;
            12'd2907: out = 16'h5A2D;
            12'd2908: out = 16'h5A25;
            12'd2909: out = 16'h5A1D;
            12'd2910: out = 16'h5A15;
            12'd2911: out = 16'h5A0E;
            12'd2912: out = 16'h5A06;
            12'd2913: out = 16'h59FE;
            12'd2914: out = 16'h59F6;
            12'd2915: out = 16'h59EE;
            12'd2916: out = 16'h59E6;
            12'd2917: out = 16'h59DE;
            12'd2918: out = 16'h59D6;
            12'd2919: out = 16'h59CE;
            12'd2920: out = 16'h59C6;
            12'd2921: out = 16'h59BF;
            12'd2922: out = 16'h59B7;
            12'd2923: out = 16'h59AF;
            12'd2924: out = 16'h59A7;
            12'd2925: out = 16'h599F;
            12'd2926: out = 16'h5997;
            12'd2927: out = 16'h5990;
            12'd2928: out = 16'h5988;
            12'd2929: out = 16'h5980;
            12'd2930: out = 16'h5978;
            12'd2931: out = 16'h5970;
            12'd2932: out = 16'h5968;
            12'd2933: out = 16'h5961;
            12'd2934: out = 16'h5959;
            12'd2935: out = 16'h5951;
            12'd2936: out = 16'h5949;
            12'd2937: out = 16'h5941;
            12'd2938: out = 16'h593A;
            12'd2939: out = 16'h5932;
            12'd2940: out = 16'h592A;
            12'd2941: out = 16'h5922;
            12'd2942: out = 16'h591B;
            12'd2943: out = 16'h5913;
            12'd2944: out = 16'h590B;
            12'd2945: out = 16'h5903;
            12'd2946: out = 16'h58FC;
            12'd2947: out = 16'h58F4;
            12'd2948: out = 16'h58EC;
            12'd2949: out = 16'h58E4;
            12'd2950: out = 16'h58DD;
            12'd2951: out = 16'h58D5;
            12'd2952: out = 16'h58CD;
            12'd2953: out = 16'h58C6;
            12'd2954: out = 16'h58BE;
            12'd2955: out = 16'h58B6;
            12'd2956: out = 16'h58AF;
            12'd2957: out = 16'h58A7;
            12'd2958: out = 16'h589F;
            12'd2959: out = 16'h5898;
            12'd2960: out = 16'h5890;
            12'd2961: out = 16'h5888;
            12'd2962: out = 16'h5881;
            12'd2963: out = 16'h5879;
            12'd2964: out = 16'h5871;
            12'd2965: out = 16'h586A;
            12'd2966: out = 16'h5862;
            12'd2967: out = 16'h585A;
            12'd2968: out = 16'h5853;
            12'd2969: out = 16'h584B;
            12'd2970: out = 16'h5844;
            12'd2971: out = 16'h583C;
            12'd2972: out = 16'h5834;
            12'd2973: out = 16'h582D;
            12'd2974: out = 16'h5825;
            12'd2975: out = 16'h581E;
            12'd2976: out = 16'h5816;
            12'd2977: out = 16'h580E;
            12'd2978: out = 16'h5807;
            12'd2979: out = 16'h57FF;
            12'd2980: out = 16'h57F8;
            12'd2981: out = 16'h57F0;
            12'd2982: out = 16'h57E9;
            12'd2983: out = 16'h57E1;
            12'd2984: out = 16'h57DA;
            12'd2985: out = 16'h57D2;
            12'd2986: out = 16'h57CB;
            12'd2987: out = 16'h57C3;
            12'd2988: out = 16'h57BB;
            12'd2989: out = 16'h57B4;
            12'd2990: out = 16'h57AC;
            12'd2991: out = 16'h57A5;
            12'd2992: out = 16'h579D;
            12'd2993: out = 16'h5796;
            12'd2994: out = 16'h578E;
            12'd2995: out = 16'h5787;
            12'd2996: out = 16'h577F;
            12'd2997: out = 16'h5778;
            12'd2998: out = 16'h5771;
            12'd2999: out = 16'h5769;
            12'd3000: out = 16'h5762;
            12'd3001: out = 16'h575A;
            12'd3002: out = 16'h5753;
            12'd3003: out = 16'h574B;
            12'd3004: out = 16'h5744;
            12'd3005: out = 16'h573C;
            12'd3006: out = 16'h5735;
            12'd3007: out = 16'h572E;
            12'd3008: out = 16'h5726;
            12'd3009: out = 16'h571F;
            12'd3010: out = 16'h5717;
            12'd3011: out = 16'h5710;
            12'd3012: out = 16'h5708;
            12'd3013: out = 16'h5701;
            12'd3014: out = 16'h56FA;
            12'd3015: out = 16'h56F2;
            12'd3016: out = 16'h56EB;
            12'd3017: out = 16'h56E4;
            12'd3018: out = 16'h56DC;
            12'd3019: out = 16'h56D5;
            12'd3020: out = 16'h56CD;
            12'd3021: out = 16'h56C6;
            12'd3022: out = 16'h56BF;
            12'd3023: out = 16'h56B7;
            12'd3024: out = 16'h56B0;
            12'd3025: out = 16'h56A9;
            12'd3026: out = 16'h56A1;
            12'd3027: out = 16'h569A;
            12'd3028: out = 16'h5693;
            12'd3029: out = 16'h568B;
            12'd3030: out = 16'h5684;
            12'd3031: out = 16'h567D;
            12'd3032: out = 16'h5676;
            12'd3033: out = 16'h566E;
            12'd3034: out = 16'h5667;
            12'd3035: out = 16'h5660;
            12'd3036: out = 16'h5658;
            12'd3037: out = 16'h5651;
            12'd3038: out = 16'h564A;
            12'd3039: out = 16'h5643;
            12'd3040: out = 16'h563B;
            12'd3041: out = 16'h5634;
            12'd3042: out = 16'h562D;
            12'd3043: out = 16'h5626;
            12'd3044: out = 16'h561E;
            12'd3045: out = 16'h5617;
            12'd3046: out = 16'h5610;
            12'd3047: out = 16'h5609;
            12'd3048: out = 16'h5601;
            12'd3049: out = 16'h55FA;
            12'd3050: out = 16'h55F3;
            12'd3051: out = 16'h55EC;
            12'd3052: out = 16'h55E4;
            12'd3053: out = 16'h55DD;
            12'd3054: out = 16'h55D6;
            12'd3055: out = 16'h55CF;
            12'd3056: out = 16'h55C8;
            12'd3057: out = 16'h55C1;
            12'd3058: out = 16'h55B9;
            12'd3059: out = 16'h55B2;
            12'd3060: out = 16'h55AB;
            12'd3061: out = 16'h55A4;
            12'd3062: out = 16'h559D;
            12'd3063: out = 16'h5596;
            12'd3064: out = 16'h558E;
            12'd3065: out = 16'h5587;
            12'd3066: out = 16'h5580;
            12'd3067: out = 16'h5579;
            12'd3068: out = 16'h5572;
            12'd3069: out = 16'h556B;
            12'd3070: out = 16'h5564;
            12'd3071: out = 16'h555C;
            12'd3072: out = 16'h5555;
            12'd3073: out = 16'h554E;
            12'd3074: out = 16'h5547;
            12'd3075: out = 16'h5540;
            12'd3076: out = 16'h5539;
            12'd3077: out = 16'h5532;
            12'd3078: out = 16'h552B;
            12'd3079: out = 16'h5524;
            12'd3080: out = 16'h551D;
            12'd3081: out = 16'h5516;
            12'd3082: out = 16'h550E;
            12'd3083: out = 16'h5507;
            12'd3084: out = 16'h5500;
            12'd3085: out = 16'h54F9;
            12'd3086: out = 16'h54F2;
            12'd3087: out = 16'h54EB;
            12'd3088: out = 16'h54E4;
            12'd3089: out = 16'h54DD;
            12'd3090: out = 16'h54D6;
            12'd3091: out = 16'h54CF;
            12'd3092: out = 16'h54C8;
            12'd3093: out = 16'h54C1;
            12'd3094: out = 16'h54BA;
            12'd3095: out = 16'h54B3;
            12'd3096: out = 16'h54AC;
            12'd3097: out = 16'h54A5;
            12'd3098: out = 16'h549E;
            12'd3099: out = 16'h5497;
            12'd3100: out = 16'h5490;
            12'd3101: out = 16'h5489;
            12'd3102: out = 16'h5482;
            12'd3103: out = 16'h547B;
            12'd3104: out = 16'h5474;
            12'd3105: out = 16'h546D;
            12'd3106: out = 16'h5466;
            12'd3107: out = 16'h545F;
            12'd3108: out = 16'h5458;
            12'd3109: out = 16'h5451;
            12'd3110: out = 16'h544A;
            12'd3111: out = 16'h5443;
            12'd3112: out = 16'h543D;
            12'd3113: out = 16'h5436;
            12'd3114: out = 16'h542F;
            12'd3115: out = 16'h5428;
            12'd3116: out = 16'h5421;
            12'd3117: out = 16'h541A;
            12'd3118: out = 16'h5413;
            12'd3119: out = 16'h540C;
            12'd3120: out = 16'h5405;
            12'd3121: out = 16'h53FE;
            12'd3122: out = 16'h53F7;
            12'd3123: out = 16'h53F1;
            12'd3124: out = 16'h53EA;
            12'd3125: out = 16'h53E3;
            12'd3126: out = 16'h53DC;
            12'd3127: out = 16'h53D5;
            12'd3128: out = 16'h53CE;
            12'd3129: out = 16'h53C7;
            12'd3130: out = 16'h53C1;
            12'd3131: out = 16'h53BA;
            12'd3132: out = 16'h53B3;
            12'd3133: out = 16'h53AC;
            12'd3134: out = 16'h53A5;
            12'd3135: out = 16'h539E;
            12'd3136: out = 16'h5398;
            12'd3137: out = 16'h5391;
            12'd3138: out = 16'h538A;
            12'd3139: out = 16'h5383;
            12'd3140: out = 16'h537C;
            12'd3141: out = 16'h5375;
            12'd3142: out = 16'h536F;
            12'd3143: out = 16'h5368;
            12'd3144: out = 16'h5361;
            12'd3145: out = 16'h535A;
            12'd3146: out = 16'h5353;
            12'd3147: out = 16'h534D;
            12'd3148: out = 16'h5346;
            12'd3149: out = 16'h533F;
            12'd3150: out = 16'h5338;
            12'd3151: out = 16'h5332;
            12'd3152: out = 16'h532B;
            12'd3153: out = 16'h5324;
            12'd3154: out = 16'h531D;
            12'd3155: out = 16'h5317;
            12'd3156: out = 16'h5310;
            12'd3157: out = 16'h5309;
            12'd3158: out = 16'h5302;
            12'd3159: out = 16'h52FC;
            12'd3160: out = 16'h52F5;
            12'd3161: out = 16'h52EE;
            12'd3162: out = 16'h52E8;
            12'd3163: out = 16'h52E1;
            12'd3164: out = 16'h52DA;
            12'd3165: out = 16'h52D3;
            12'd3166: out = 16'h52CD;
            12'd3167: out = 16'h52C6;
            12'd3168: out = 16'h52BF;
            12'd3169: out = 16'h52B9;
            12'd3170: out = 16'h52B2;
            12'd3171: out = 16'h52AB;
            12'd3172: out = 16'h52A5;
            12'd3173: out = 16'h529E;
            12'd3174: out = 16'h5297;
            12'd3175: out = 16'h5291;
            12'd3176: out = 16'h528A;
            12'd3177: out = 16'h5283;
            12'd3178: out = 16'h527D;
            12'd3179: out = 16'h5276;
            12'd3180: out = 16'h526F;
            12'd3181: out = 16'h5269;
            12'd3182: out = 16'h5262;
            12'd3183: out = 16'h525C;
            12'd3184: out = 16'h5255;
            12'd3185: out = 16'h524E;
            12'd3186: out = 16'h5248;
            12'd3187: out = 16'h5241;
            12'd3188: out = 16'h523A;
            12'd3189: out = 16'h5234;
            12'd3190: out = 16'h522D;
            12'd3191: out = 16'h5227;
            12'd3192: out = 16'h5220;
            12'd3193: out = 16'h5219;
            12'd3194: out = 16'h5213;
            12'd3195: out = 16'h520C;
            12'd3196: out = 16'h5206;
            12'd3197: out = 16'h51FF;
            12'd3198: out = 16'h51F9;
            12'd3199: out = 16'h51F2;
            12'd3200: out = 16'h51EC;
            12'd3201: out = 16'h51E5;
            12'd3202: out = 16'h51DE;
            12'd3203: out = 16'h51D8;
            12'd3204: out = 16'h51D1;
            12'd3205: out = 16'h51CB;
            12'd3206: out = 16'h51C4;
            12'd3207: out = 16'h51BE;
            12'd3208: out = 16'h51B7;
            12'd3209: out = 16'h51B1;
            12'd3210: out = 16'h51AA;
            12'd3211: out = 16'h51A4;
            12'd3212: out = 16'h519D;
            12'd3213: out = 16'h5197;
            12'd3214: out = 16'h5190;
            12'd3215: out = 16'h518A;
            12'd3216: out = 16'h5183;
            12'd3217: out = 16'h517D;
            12'd3218: out = 16'h5176;
            12'd3219: out = 16'h5170;
            12'd3220: out = 16'h5169;
            12'd3221: out = 16'h5163;
            12'd3222: out = 16'h515C;
            12'd3223: out = 16'h5156;
            12'd3224: out = 16'h514F;
            12'd3225: out = 16'h5149;
            12'd3226: out = 16'h5142;
            12'd3227: out = 16'h513C;
            12'd3228: out = 16'h5136;
            12'd3229: out = 16'h512F;
            12'd3230: out = 16'h5129;
            12'd3231: out = 16'h5122;
            12'd3232: out = 16'h511C;
            12'd3233: out = 16'h5115;
            12'd3234: out = 16'h510F;
            12'd3235: out = 16'h5109;
            12'd3236: out = 16'h5102;
            12'd3237: out = 16'h50FC;
            12'd3238: out = 16'h50F5;
            12'd3239: out = 16'h50EF;
            12'd3240: out = 16'h50E9;
            12'd3241: out = 16'h50E2;
            12'd3242: out = 16'h50DC;
            12'd3243: out = 16'h50D5;
            12'd3244: out = 16'h50CF;
            12'd3245: out = 16'h50C9;
            12'd3246: out = 16'h50C2;
            12'd3247: out = 16'h50BC;
            12'd3248: out = 16'h50B6;
            12'd3249: out = 16'h50AF;
            12'd3250: out = 16'h50A9;
            12'd3251: out = 16'h50A3;
            12'd3252: out = 16'h509C;
            12'd3253: out = 16'h5096;
            12'd3254: out = 16'h508F;
            12'd3255: out = 16'h5089;
            12'd3256: out = 16'h5083;
            12'd3257: out = 16'h507D;
            12'd3258: out = 16'h5076;
            12'd3259: out = 16'h5070;
            12'd3260: out = 16'h506A;
            12'd3261: out = 16'h5063;
            12'd3262: out = 16'h505D;
            12'd3263: out = 16'h5057;
            12'd3264: out = 16'h5050;
            12'd3265: out = 16'h504A;
            12'd3266: out = 16'h5044;
            12'd3267: out = 16'h503D;
            12'd3268: out = 16'h5037;
            12'd3269: out = 16'h5031;
            12'd3270: out = 16'h502B;
            12'd3271: out = 16'h5024;
            12'd3272: out = 16'h501E;
            12'd3273: out = 16'h5018;
            12'd3274: out = 16'h5012;
            12'd3275: out = 16'h500B;
            12'd3276: out = 16'h5005;
            12'd3277: out = 16'h4FFF;
            12'd3278: out = 16'h4FF9;
            12'd3279: out = 16'h4FF2;
            12'd3280: out = 16'h4FEC;
            12'd3281: out = 16'h4FE6;
            12'd3282: out = 16'h4FE0;
            12'd3283: out = 16'h4FD9;
            12'd3284: out = 16'h4FD3;
            12'd3285: out = 16'h4FCD;
            12'd3286: out = 16'h4FC7;
            12'd3287: out = 16'h4FC0;
            12'd3288: out = 16'h4FBA;
            12'd3289: out = 16'h4FB4;
            12'd3290: out = 16'h4FAE;
            12'd3291: out = 16'h4FA8;
            12'd3292: out = 16'h4FA1;
            12'd3293: out = 16'h4F9B;
            12'd3294: out = 16'h4F95;
            12'd3295: out = 16'h4F8F;
            12'd3296: out = 16'h4F89;
            12'd3297: out = 16'h4F83;
            12'd3298: out = 16'h4F7C;
            12'd3299: out = 16'h4F76;
            12'd3300: out = 16'h4F70;
            12'd3301: out = 16'h4F6A;
            12'd3302: out = 16'h4F64;
            12'd3303: out = 16'h4F5E;
            12'd3304: out = 16'h4F57;
            12'd3305: out = 16'h4F51;
            12'd3306: out = 16'h4F4B;
            12'd3307: out = 16'h4F45;
            12'd3308: out = 16'h4F3F;
            12'd3309: out = 16'h4F39;
            12'd3310: out = 16'h4F33;
            12'd3311: out = 16'h4F2C;
            12'd3312: out = 16'h4F26;
            12'd3313: out = 16'h4F20;
            12'd3314: out = 16'h4F1A;
            12'd3315: out = 16'h4F14;
            12'd3316: out = 16'h4F0E;
            12'd3317: out = 16'h4F08;
            12'd3318: out = 16'h4F02;
            12'd3319: out = 16'h4EFC;
            12'd3320: out = 16'h4EF6;
            12'd3321: out = 16'h4EEF;
            12'd3322: out = 16'h4EE9;
            12'd3323: out = 16'h4EE3;
            12'd3324: out = 16'h4EDD;
            12'd3325: out = 16'h4ED7;
            12'd3326: out = 16'h4ED1;
            12'd3327: out = 16'h4ECB;
            12'd3328: out = 16'h4EC5;
            12'd3329: out = 16'h4EBF;
            12'd3330: out = 16'h4EB9;
            12'd3331: out = 16'h4EB3;
            12'd3332: out = 16'h4EAD;
            12'd3333: out = 16'h4EA7;
            12'd3334: out = 16'h4EA1;
            12'd3335: out = 16'h4E9B;
            12'd3336: out = 16'h4E95;
            12'd3337: out = 16'h4E8F;
            12'd3338: out = 16'h4E89;
            12'd3339: out = 16'h4E82;
            12'd3340: out = 16'h4E7C;
            12'd3341: out = 16'h4E76;
            12'd3342: out = 16'h4E70;
            12'd3343: out = 16'h4E6A;
            12'd3344: out = 16'h4E64;
            12'd3345: out = 16'h4E5E;
            12'd3346: out = 16'h4E58;
            12'd3347: out = 16'h4E52;
            12'd3348: out = 16'h4E4C;
            12'd3349: out = 16'h4E46;
            12'd3350: out = 16'h4E40;
            12'd3351: out = 16'h4E3B;
            12'd3352: out = 16'h4E35;
            12'd3353: out = 16'h4E2F;
            12'd3354: out = 16'h4E29;
            12'd3355: out = 16'h4E23;
            12'd3356: out = 16'h4E1D;
            12'd3357: out = 16'h4E17;
            12'd3358: out = 16'h4E11;
            12'd3359: out = 16'h4E0B;
            12'd3360: out = 16'h4E05;
            12'd3361: out = 16'h4DFF;
            12'd3362: out = 16'h4DF9;
            12'd3363: out = 16'h4DF3;
            12'd3364: out = 16'h4DED;
            12'd3365: out = 16'h4DE7;
            12'd3366: out = 16'h4DE1;
            12'd3367: out = 16'h4DDB;
            12'd3368: out = 16'h4DD5;
            12'd3369: out = 16'h4DD0;
            12'd3370: out = 16'h4DCA;
            12'd3371: out = 16'h4DC4;
            12'd3372: out = 16'h4DBE;
            12'd3373: out = 16'h4DB8;
            12'd3374: out = 16'h4DB2;
            12'd3375: out = 16'h4DAC;
            12'd3376: out = 16'h4DA6;
            12'd3377: out = 16'h4DA0;
            12'd3378: out = 16'h4D9A;
            12'd3379: out = 16'h4D95;
            12'd3380: out = 16'h4D8F;
            12'd3381: out = 16'h4D89;
            12'd3382: out = 16'h4D83;
            12'd3383: out = 16'h4D7D;
            12'd3384: out = 16'h4D77;
            12'd3385: out = 16'h4D71;
            12'd3386: out = 16'h4D6C;
            12'd3387: out = 16'h4D66;
            12'd3388: out = 16'h4D60;
            12'd3389: out = 16'h4D5A;
            12'd3390: out = 16'h4D54;
            12'd3391: out = 16'h4D4E;
            12'd3392: out = 16'h4D48;
            12'd3393: out = 16'h4D43;
            12'd3394: out = 16'h4D3D;
            12'd3395: out = 16'h4D37;
            12'd3396: out = 16'h4D31;
            12'd3397: out = 16'h4D2B;
            12'd3398: out = 16'h4D26;
            12'd3399: out = 16'h4D20;
            12'd3400: out = 16'h4D1A;
            12'd3401: out = 16'h4D14;
            12'd3402: out = 16'h4D0E;
            12'd3403: out = 16'h4D09;
            12'd3404: out = 16'h4D03;
            12'd3405: out = 16'h4CFD;
            12'd3406: out = 16'h4CF7;
            12'd3407: out = 16'h4CF1;
            12'd3408: out = 16'h4CEC;
            12'd3409: out = 16'h4CE6;
            12'd3410: out = 16'h4CE0;
            12'd3411: out = 16'h4CDA;
            12'd3412: out = 16'h4CD4;
            12'd3413: out = 16'h4CCF;
            12'd3414: out = 16'h4CC9;
            12'd3415: out = 16'h4CC3;
            12'd3416: out = 16'h4CBD;
            12'd3417: out = 16'h4CB8;
            12'd3418: out = 16'h4CB2;
            12'd3419: out = 16'h4CAC;
            12'd3420: out = 16'h4CA6;
            12'd3421: out = 16'h4CA1;
            12'd3422: out = 16'h4C9B;
            12'd3423: out = 16'h4C95;
            12'd3424: out = 16'h4C90;
            12'd3425: out = 16'h4C8A;
            12'd3426: out = 16'h4C84;
            12'd3427: out = 16'h4C7E;
            12'd3428: out = 16'h4C79;
            12'd3429: out = 16'h4C73;
            12'd3430: out = 16'h4C6D;
            12'd3431: out = 16'h4C68;
            12'd3432: out = 16'h4C62;
            12'd3433: out = 16'h4C5C;
            12'd3434: out = 16'h4C56;
            12'd3435: out = 16'h4C51;
            12'd3436: out = 16'h4C4B;
            12'd3437: out = 16'h4C45;
            12'd3438: out = 16'h4C40;
            12'd3439: out = 16'h4C3A;
            12'd3440: out = 16'h4C34;
            12'd3441: out = 16'h4C2F;
            12'd3442: out = 16'h4C29;
            12'd3443: out = 16'h4C23;
            12'd3444: out = 16'h4C1E;
            12'd3445: out = 16'h4C18;
            12'd3446: out = 16'h4C12;
            12'd3447: out = 16'h4C0D;
            12'd3448: out = 16'h4C07;
            12'd3449: out = 16'h4C01;
            12'd3450: out = 16'h4BFC;
            12'd3451: out = 16'h4BF6;
            12'd3452: out = 16'h4BF1;
            12'd3453: out = 16'h4BEB;
            12'd3454: out = 16'h4BE5;
            12'd3455: out = 16'h4BE0;
            12'd3456: out = 16'h4BDA;
            12'd3457: out = 16'h4BD4;
            12'd3458: out = 16'h4BCF;
            12'd3459: out = 16'h4BC9;
            12'd3460: out = 16'h4BC4;
            12'd3461: out = 16'h4BBE;
            12'd3462: out = 16'h4BB8;
            12'd3463: out = 16'h4BB3;
            12'd3464: out = 16'h4BAD;
            12'd3465: out = 16'h4BA8;
            12'd3466: out = 16'h4BA2;
            12'd3467: out = 16'h4B9C;
            12'd3468: out = 16'h4B97;
            12'd3469: out = 16'h4B91;
            12'd3470: out = 16'h4B8C;
            12'd3471: out = 16'h4B86;
            12'd3472: out = 16'h4B81;
            12'd3473: out = 16'h4B7B;
            12'd3474: out = 16'h4B75;
            12'd3475: out = 16'h4B70;
            12'd3476: out = 16'h4B6A;
            12'd3477: out = 16'h4B65;
            12'd3478: out = 16'h4B5F;
            12'd3479: out = 16'h4B5A;
            12'd3480: out = 16'h4B54;
            12'd3481: out = 16'h4B4F;
            12'd3482: out = 16'h4B49;
            12'd3483: out = 16'h4B44;
            12'd3484: out = 16'h4B3E;
            12'd3485: out = 16'h4B38;
            12'd3486: out = 16'h4B33;
            12'd3487: out = 16'h4B2D;
            12'd3488: out = 16'h4B28;
            12'd3489: out = 16'h4B22;
            12'd3490: out = 16'h4B1D;
            12'd3491: out = 16'h4B17;
            12'd3492: out = 16'h4B12;
            12'd3493: out = 16'h4B0C;
            12'd3494: out = 16'h4B07;
            12'd3495: out = 16'h4B01;
            12'd3496: out = 16'h4AFC;
            12'd3497: out = 16'h4AF6;
            12'd3498: out = 16'h4AF1;
            12'd3499: out = 16'h4AEB;
            12'd3500: out = 16'h4AE6;
            12'd3501: out = 16'h4AE0;
            12'd3502: out = 16'h4ADB;
            12'd3503: out = 16'h4AD6;
            12'd3504: out = 16'h4AD0;
            12'd3505: out = 16'h4ACB;
            12'd3506: out = 16'h4AC5;
            12'd3507: out = 16'h4AC0;
            12'd3508: out = 16'h4ABA;
            12'd3509: out = 16'h4AB5;
            12'd3510: out = 16'h4AAF;
            12'd3511: out = 16'h4AAA;
            12'd3512: out = 16'h4AA4;
            12'd3513: out = 16'h4A9F;
            12'd3514: out = 16'h4A9A;
            12'd3515: out = 16'h4A94;
            12'd3516: out = 16'h4A8F;
            12'd3517: out = 16'h4A89;
            12'd3518: out = 16'h4A84;
            12'd3519: out = 16'h4A7E;
            12'd3520: out = 16'h4A79;
            12'd3521: out = 16'h4A74;
            12'd3522: out = 16'h4A6E;
            12'd3523: out = 16'h4A69;
            12'd3524: out = 16'h4A63;
            12'd3525: out = 16'h4A5E;
            12'd3526: out = 16'h4A59;
            12'd3527: out = 16'h4A53;
            12'd3528: out = 16'h4A4E;
            12'd3529: out = 16'h4A48;
            12'd3530: out = 16'h4A43;
            12'd3531: out = 16'h4A3E;
            12'd3532: out = 16'h4A38;
            12'd3533: out = 16'h4A33;
            12'd3534: out = 16'h4A2D;
            12'd3535: out = 16'h4A28;
            12'd3536: out = 16'h4A23;
            12'd3537: out = 16'h4A1D;
            12'd3538: out = 16'h4A18;
            12'd3539: out = 16'h4A13;
            12'd3540: out = 16'h4A0D;
            12'd3541: out = 16'h4A08;
            12'd3542: out = 16'h4A03;
            12'd3543: out = 16'h49FD;
            12'd3544: out = 16'h49F8;
            12'd3545: out = 16'h49F3;
            12'd3546: out = 16'h49ED;
            12'd3547: out = 16'h49E8;
            12'd3548: out = 16'h49E3;
            12'd3549: out = 16'h49DD;
            12'd3550: out = 16'h49D8;
            12'd3551: out = 16'h49D3;
            12'd3552: out = 16'h49CD;
            12'd3553: out = 16'h49C8;
            12'd3554: out = 16'h49C3;
            12'd3555: out = 16'h49BD;
            12'd3556: out = 16'h49B8;
            12'd3557: out = 16'h49B3;
            12'd3558: out = 16'h49AD;
            12'd3559: out = 16'h49A8;
            12'd3560: out = 16'h49A3;
            12'd3561: out = 16'h499E;
            12'd3562: out = 16'h4998;
            12'd3563: out = 16'h4993;
            12'd3564: out = 16'h498E;
            12'd3565: out = 16'h4988;
            12'd3566: out = 16'h4983;
            12'd3567: out = 16'h497E;
            12'd3568: out = 16'h4979;
            12'd3569: out = 16'h4973;
            12'd3570: out = 16'h496E;
            12'd3571: out = 16'h4969;
            12'd3572: out = 16'h4963;
            12'd3573: out = 16'h495E;
            12'd3574: out = 16'h4959;
            12'd3575: out = 16'h4954;
            12'd3576: out = 16'h494E;
            12'd3577: out = 16'h4949;
            12'd3578: out = 16'h4944;
            12'd3579: out = 16'h493F;
            12'd3580: out = 16'h4939;
            12'd3581: out = 16'h4934;
            12'd3582: out = 16'h492F;
            12'd3583: out = 16'h492A;
            12'd3584: out = 16'h4925;
            12'd3585: out = 16'h491F;
            12'd3586: out = 16'h491A;
            12'd3587: out = 16'h4915;
            12'd3588: out = 16'h4910;
            12'd3589: out = 16'h490A;
            12'd3590: out = 16'h4905;
            12'd3591: out = 16'h4900;
            12'd3592: out = 16'h48FB;
            12'd3593: out = 16'h48F6;
            12'd3594: out = 16'h48F0;
            12'd3595: out = 16'h48EB;
            12'd3596: out = 16'h48E6;
            12'd3597: out = 16'h48E1;
            12'd3598: out = 16'h48DC;
            12'd3599: out = 16'h48D7;
            12'd3600: out = 16'h48D1;
            12'd3601: out = 16'h48CC;
            12'd3602: out = 16'h48C7;
            12'd3603: out = 16'h48C2;
            12'd3604: out = 16'h48BD;
            12'd3605: out = 16'h48B7;
            12'd3606: out = 16'h48B2;
            12'd3607: out = 16'h48AD;
            12'd3608: out = 16'h48A8;
            12'd3609: out = 16'h48A3;
            12'd3610: out = 16'h489E;
            12'd3611: out = 16'h4899;
            12'd3612: out = 16'h4893;
            12'd3613: out = 16'h488E;
            12'd3614: out = 16'h4889;
            12'd3615: out = 16'h4884;
            12'd3616: out = 16'h487F;
            12'd3617: out = 16'h487A;
            12'd3618: out = 16'h4875;
            12'd3619: out = 16'h486F;
            12'd3620: out = 16'h486A;
            12'd3621: out = 16'h4865;
            12'd3622: out = 16'h4860;
            12'd3623: out = 16'h485B;
            12'd3624: out = 16'h4856;
            12'd3625: out = 16'h4851;
            12'd3626: out = 16'h484C;
            12'd3627: out = 16'h4847;
            12'd3628: out = 16'h4841;
            12'd3629: out = 16'h483C;
            12'd3630: out = 16'h4837;
            12'd3631: out = 16'h4832;
            12'd3632: out = 16'h482D;
            12'd3633: out = 16'h4828;
            12'd3634: out = 16'h4823;
            12'd3635: out = 16'h481E;
            12'd3636: out = 16'h4819;
            12'd3637: out = 16'h4814;
            12'd3638: out = 16'h480F;
            12'd3639: out = 16'h480A;
            12'd3640: out = 16'h4805;
            12'd3641: out = 16'h47FF;
            12'd3642: out = 16'h47FA;
            12'd3643: out = 16'h47F5;
            12'd3644: out = 16'h47F0;
            12'd3645: out = 16'h47EB;
            12'd3646: out = 16'h47E6;
            12'd3647: out = 16'h47E1;
            12'd3648: out = 16'h47DC;
            12'd3649: out = 16'h47D7;
            12'd3650: out = 16'h47D2;
            12'd3651: out = 16'h47CD;
            12'd3652: out = 16'h47C8;
            12'd3653: out = 16'h47C3;
            12'd3654: out = 16'h47BE;
            12'd3655: out = 16'h47B9;
            12'd3656: out = 16'h47B4;
            12'd3657: out = 16'h47AF;
            12'd3658: out = 16'h47AA;
            12'd3659: out = 16'h47A5;
            12'd3660: out = 16'h47A0;
            12'd3661: out = 16'h479B;
            12'd3662: out = 16'h4796;
            12'd3663: out = 16'h4791;
            12'd3664: out = 16'h478C;
            12'd3665: out = 16'h4787;
            12'd3666: out = 16'h4782;
            12'd3667: out = 16'h477D;
            12'd3668: out = 16'h4778;
            12'd3669: out = 16'h4773;
            12'd3670: out = 16'h476E;
            12'd3671: out = 16'h4769;
            12'd3672: out = 16'h4764;
            12'd3673: out = 16'h475F;
            12'd3674: out = 16'h475A;
            12'd3675: out = 16'h4755;
            12'd3676: out = 16'h4750;
            12'd3677: out = 16'h474B;
            12'd3678: out = 16'h4746;
            12'd3679: out = 16'h4741;
            12'd3680: out = 16'h473C;
            12'd3681: out = 16'h4737;
            12'd3682: out = 16'h4732;
            12'd3683: out = 16'h472D;
            12'd3684: out = 16'h4728;
            12'd3685: out = 16'h4723;
            12'd3686: out = 16'h471E;
            12'd3687: out = 16'h4719;
            12'd3688: out = 16'h4715;
            12'd3689: out = 16'h4710;
            12'd3690: out = 16'h470B;
            12'd3691: out = 16'h4706;
            12'd3692: out = 16'h4701;
            12'd3693: out = 16'h46FC;
            12'd3694: out = 16'h46F7;
            12'd3695: out = 16'h46F2;
            12'd3696: out = 16'h46ED;
            12'd3697: out = 16'h46E8;
            12'd3698: out = 16'h46E3;
            12'd3699: out = 16'h46DE;
            12'd3700: out = 16'h46DA;
            12'd3701: out = 16'h46D5;
            12'd3702: out = 16'h46D0;
            12'd3703: out = 16'h46CB;
            12'd3704: out = 16'h46C6;
            12'd3705: out = 16'h46C1;
            12'd3706: out = 16'h46BC;
            12'd3707: out = 16'h46B7;
            12'd3708: out = 16'h46B2;
            12'd3709: out = 16'h46AE;
            12'd3710: out = 16'h46A9;
            12'd3711: out = 16'h46A4;
            12'd3712: out = 16'h469F;
            12'd3713: out = 16'h469A;
            12'd3714: out = 16'h4695;
            12'd3715: out = 16'h4690;
            12'd3716: out = 16'h468B;
            12'd3717: out = 16'h4687;
            12'd3718: out = 16'h4682;
            12'd3719: out = 16'h467D;
            12'd3720: out = 16'h4678;
            12'd3721: out = 16'h4673;
            12'd3722: out = 16'h466E;
            12'd3723: out = 16'h4669;
            12'd3724: out = 16'h4665;
            12'd3725: out = 16'h4660;
            12'd3726: out = 16'h465B;
            12'd3727: out = 16'h4656;
            12'd3728: out = 16'h4651;
            12'd3729: out = 16'h464C;
            12'd3730: out = 16'h4648;
            12'd3731: out = 16'h4643;
            12'd3732: out = 16'h463E;
            12'd3733: out = 16'h4639;
            12'd3734: out = 16'h4634;
            12'd3735: out = 16'h4630;
            12'd3736: out = 16'h462B;
            12'd3737: out = 16'h4626;
            12'd3738: out = 16'h4621;
            12'd3739: out = 16'h461C;
            12'd3740: out = 16'h4618;
            12'd3741: out = 16'h4613;
            12'd3742: out = 16'h460E;
            12'd3743: out = 16'h4609;
            12'd3744: out = 16'h4604;
            12'd3745: out = 16'h4600;
            12'd3746: out = 16'h45FB;
            12'd3747: out = 16'h45F6;
            12'd3748: out = 16'h45F1;
            12'd3749: out = 16'h45EC;
            12'd3750: out = 16'h45E8;
            12'd3751: out = 16'h45E3;
            12'd3752: out = 16'h45DE;
            12'd3753: out = 16'h45D9;
            12'd3754: out = 16'h45D5;
            12'd3755: out = 16'h45D0;
            12'd3756: out = 16'h45CB;
            12'd3757: out = 16'h45C6;
            12'd3758: out = 16'h45C2;
            12'd3759: out = 16'h45BD;
            12'd3760: out = 16'h45B8;
            12'd3761: out = 16'h45B3;
            12'd3762: out = 16'h45AF;
            12'd3763: out = 16'h45AA;
            12'd3764: out = 16'h45A5;
            12'd3765: out = 16'h45A0;
            12'd3766: out = 16'h459C;
            12'd3767: out = 16'h4597;
            12'd3768: out = 16'h4592;
            12'd3769: out = 16'h458D;
            12'd3770: out = 16'h4589;
            12'd3771: out = 16'h4584;
            12'd3772: out = 16'h457F;
            12'd3773: out = 16'h457B;
            12'd3774: out = 16'h4576;
            12'd3775: out = 16'h4571;
            12'd3776: out = 16'h456C;
            12'd3777: out = 16'h4568;
            12'd3778: out = 16'h4563;
            12'd3779: out = 16'h455E;
            12'd3780: out = 16'h455A;
            12'd3781: out = 16'h4555;
            12'd3782: out = 16'h4550;
            12'd3783: out = 16'h454C;
            12'd3784: out = 16'h4547;
            12'd3785: out = 16'h4542;
            12'd3786: out = 16'h453E;
            12'd3787: out = 16'h4539;
            12'd3788: out = 16'h4534;
            12'd3789: out = 16'h452F;
            12'd3790: out = 16'h452B;
            12'd3791: out = 16'h4526;
            12'd3792: out = 16'h4521;
            12'd3793: out = 16'h451D;
            12'd3794: out = 16'h4518;
            12'd3795: out = 16'h4513;
            12'd3796: out = 16'h450F;
            12'd3797: out = 16'h450A;
            12'd3798: out = 16'h4506;
            12'd3799: out = 16'h4501;
            12'd3800: out = 16'h44FC;
            12'd3801: out = 16'h44F8;
            12'd3802: out = 16'h44F3;
            12'd3803: out = 16'h44EE;
            12'd3804: out = 16'h44EA;
            12'd3805: out = 16'h44E5;
            12'd3806: out = 16'h44E0;
            12'd3807: out = 16'h44DC;
            12'd3808: out = 16'h44D7;
            12'd3809: out = 16'h44D2;
            12'd3810: out = 16'h44CE;
            12'd3811: out = 16'h44C9;
            12'd3812: out = 16'h44C5;
            12'd3813: out = 16'h44C0;
            12'd3814: out = 16'h44BB;
            12'd3815: out = 16'h44B7;
            12'd3816: out = 16'h44B2;
            12'd3817: out = 16'h44AE;
            12'd3818: out = 16'h44A9;
            12'd3819: out = 16'h44A4;
            12'd3820: out = 16'h44A0;
            12'd3821: out = 16'h449B;
            12'd3822: out = 16'h4497;
            12'd3823: out = 16'h4492;
            12'd3824: out = 16'h448D;
            12'd3825: out = 16'h4489;
            12'd3826: out = 16'h4484;
            12'd3827: out = 16'h4480;
            12'd3828: out = 16'h447B;
            12'd3829: out = 16'h4476;
            12'd3830: out = 16'h4472;
            12'd3831: out = 16'h446D;
            12'd3832: out = 16'h4469;
            12'd3833: out = 16'h4464;
            12'd3834: out = 16'h4460;
            12'd3835: out = 16'h445B;
            12'd3836: out = 16'h4456;
            12'd3837: out = 16'h4452;
            12'd3838: out = 16'h444D;
            12'd3839: out = 16'h4449;
            12'd3840: out = 16'h4444;
            12'd3841: out = 16'h4440;
            12'd3842: out = 16'h443B;
            12'd3843: out = 16'h4437;
            12'd3844: out = 16'h4432;
            12'd3845: out = 16'h442E;
            12'd3846: out = 16'h4429;
            12'd3847: out = 16'h4424;
            12'd3848: out = 16'h4420;
            12'd3849: out = 16'h441B;
            12'd3850: out = 16'h4417;
            12'd3851: out = 16'h4412;
            12'd3852: out = 16'h440E;
            12'd3853: out = 16'h4409;
            12'd3854: out = 16'h4405;
            12'd3855: out = 16'h4400;
            12'd3856: out = 16'h43FC;
            12'd3857: out = 16'h43F7;
            12'd3858: out = 16'h43F3;
            12'd3859: out = 16'h43EE;
            12'd3860: out = 16'h43EA;
            12'd3861: out = 16'h43E5;
            12'd3862: out = 16'h43E1;
            12'd3863: out = 16'h43DC;
            12'd3864: out = 16'h43D8;
            12'd3865: out = 16'h43D3;
            12'd3866: out = 16'h43CF;
            12'd3867: out = 16'h43CA;
            12'd3868: out = 16'h43C6;
            12'd3869: out = 16'h43C1;
            12'd3870: out = 16'h43BD;
            12'd3871: out = 16'h43B8;
            12'd3872: out = 16'h43B4;
            12'd3873: out = 16'h43AF;
            12'd3874: out = 16'h43AB;
            12'd3875: out = 16'h43A6;
            12'd3876: out = 16'h43A2;
            12'd3877: out = 16'h439D;
            12'd3878: out = 16'h4399;
            12'd3879: out = 16'h4395;
            12'd3880: out = 16'h4390;
            12'd3881: out = 16'h438C;
            12'd3882: out = 16'h4387;
            12'd3883: out = 16'h4383;
            12'd3884: out = 16'h437E;
            12'd3885: out = 16'h437A;
            12'd3886: out = 16'h4375;
            12'd3887: out = 16'h4371;
            12'd3888: out = 16'h436D;
            12'd3889: out = 16'h4368;
            12'd3890: out = 16'h4364;
            12'd3891: out = 16'h435F;
            12'd3892: out = 16'h435B;
            12'd3893: out = 16'h4356;
            12'd3894: out = 16'h4352;
            12'd3895: out = 16'h434D;
            12'd3896: out = 16'h4349;
            12'd3897: out = 16'h4345;
            12'd3898: out = 16'h4340;
            12'd3899: out = 16'h433C;
            12'd3900: out = 16'h4337;
            12'd3901: out = 16'h4333;
            12'd3902: out = 16'h432F;
            12'd3903: out = 16'h432A;
            12'd3904: out = 16'h4326;
            12'd3905: out = 16'h4321;
            12'd3906: out = 16'h431D;
            12'd3907: out = 16'h4319;
            12'd3908: out = 16'h4314;
            12'd3909: out = 16'h4310;
            12'd3910: out = 16'h430B;
            12'd3911: out = 16'h4307;
            12'd3912: out = 16'h4303;
            12'd3913: out = 16'h42FE;
            12'd3914: out = 16'h42FA;
            12'd3915: out = 16'h42F5;
            12'd3916: out = 16'h42F1;
            12'd3917: out = 16'h42ED;
            12'd3918: out = 16'h42E8;
            12'd3919: out = 16'h42E4;
            12'd3920: out = 16'h42E0;
            12'd3921: out = 16'h42DB;
            12'd3922: out = 16'h42D7;
            12'd3923: out = 16'h42D3;
            12'd3924: out = 16'h42CE;
            12'd3925: out = 16'h42CA;
            12'd3926: out = 16'h42C5;
            12'd3927: out = 16'h42C1;
            12'd3928: out = 16'h42BD;
            12'd3929: out = 16'h42B8;
            12'd3930: out = 16'h42B4;
            12'd3931: out = 16'h42B0;
            12'd3932: out = 16'h42AB;
            12'd3933: out = 16'h42A7;
            12'd3934: out = 16'h42A3;
            12'd3935: out = 16'h429E;
            12'd3936: out = 16'h429A;
            12'd3937: out = 16'h4296;
            12'd3938: out = 16'h4291;
            12'd3939: out = 16'h428D;
            12'd3940: out = 16'h4289;
            12'd3941: out = 16'h4284;
            12'd3942: out = 16'h4280;
            12'd3943: out = 16'h427C;
            12'd3944: out = 16'h4277;
            12'd3945: out = 16'h4273;
            12'd3946: out = 16'h426F;
            12'd3947: out = 16'h426A;
            12'd3948: out = 16'h4266;
            12'd3949: out = 16'h4262;
            12'd3950: out = 16'h425E;
            12'd3951: out = 16'h4259;
            12'd3952: out = 16'h4255;
            12'd3953: out = 16'h4251;
            12'd3954: out = 16'h424C;
            12'd3955: out = 16'h4248;
            12'd3956: out = 16'h4244;
            12'd3957: out = 16'h4240;
            12'd3958: out = 16'h423B;
            12'd3959: out = 16'h4237;
            12'd3960: out = 16'h4233;
            12'd3961: out = 16'h422E;
            12'd3962: out = 16'h422A;
            12'd3963: out = 16'h4226;
            12'd3964: out = 16'h4222;
            12'd3965: out = 16'h421D;
            12'd3966: out = 16'h4219;
            12'd3967: out = 16'h4215;
            12'd3968: out = 16'h4211;
            12'd3969: out = 16'h420C;
            12'd3970: out = 16'h4208;
            12'd3971: out = 16'h4204;
            12'd3972: out = 16'h41FF;
            12'd3973: out = 16'h41FB;
            12'd3974: out = 16'h41F7;
            12'd3975: out = 16'h41F3;
            12'd3976: out = 16'h41EE;
            12'd3977: out = 16'h41EA;
            12'd3978: out = 16'h41E6;
            12'd3979: out = 16'h41E2;
            12'd3980: out = 16'h41DE;
            12'd3981: out = 16'h41D9;
            12'd3982: out = 16'h41D5;
            12'd3983: out = 16'h41D1;
            12'd3984: out = 16'h41CD;
            12'd3985: out = 16'h41C8;
            12'd3986: out = 16'h41C4;
            12'd3987: out = 16'h41C0;
            12'd3988: out = 16'h41BC;
            12'd3989: out = 16'h41B7;
            12'd3990: out = 16'h41B3;
            12'd3991: out = 16'h41AF;
            12'd3992: out = 16'h41AB;
            12'd3993: out = 16'h41A7;
            12'd3994: out = 16'h41A2;
            12'd3995: out = 16'h419E;
            12'd3996: out = 16'h419A;
            12'd3997: out = 16'h4196;
            12'd3998: out = 16'h4192;
            12'd3999: out = 16'h418D;
            12'd4000: out = 16'h4189;
            12'd4001: out = 16'h4185;
            12'd4002: out = 16'h4181;
            12'd4003: out = 16'h417D;
            12'd4004: out = 16'h4178;
            12'd4005: out = 16'h4174;
            12'd4006: out = 16'h4170;
            12'd4007: out = 16'h416C;
            12'd4008: out = 16'h4168;
            12'd4009: out = 16'h4164;
            12'd4010: out = 16'h415F;
            12'd4011: out = 16'h415B;
            12'd4012: out = 16'h4157;
            12'd4013: out = 16'h4153;
            12'd4014: out = 16'h414F;
            12'd4015: out = 16'h414B;
            12'd4016: out = 16'h4146;
            12'd4017: out = 16'h4142;
            12'd4018: out = 16'h413E;
            12'd4019: out = 16'h413A;
            12'd4020: out = 16'h4136;
            12'd4021: out = 16'h4132;
            12'd4022: out = 16'h412D;
            12'd4023: out = 16'h4129;
            12'd4024: out = 16'h4125;
            12'd4025: out = 16'h4121;
            12'd4026: out = 16'h411D;
            12'd4027: out = 16'h4119;
            12'd4028: out = 16'h4115;
            12'd4029: out = 16'h4110;
            12'd4030: out = 16'h410C;
            12'd4031: out = 16'h4108;
            12'd4032: out = 16'h4104;
            12'd4033: out = 16'h4100;
            12'd4034: out = 16'h40FC;
            12'd4035: out = 16'h40F8;
            12'd4036: out = 16'h40F4;
            12'd4037: out = 16'h40EF;
            12'd4038: out = 16'h40EB;
            12'd4039: out = 16'h40E7;
            12'd4040: out = 16'h40E3;
            12'd4041: out = 16'h40DF;
            12'd4042: out = 16'h40DB;
            12'd4043: out = 16'h40D7;
            12'd4044: out = 16'h40D3;
            12'd4045: out = 16'h40CF;
            12'd4046: out = 16'h40CA;
            12'd4047: out = 16'h40C6;
            12'd4048: out = 16'h40C2;
            12'd4049: out = 16'h40BE;
            12'd4050: out = 16'h40BA;
            12'd4051: out = 16'h40B6;
            12'd4052: out = 16'h40B2;
            12'd4053: out = 16'h40AE;
            12'd4054: out = 16'h40AA;
            12'd4055: out = 16'h40A6;
            12'd4056: out = 16'h40A2;
            12'd4057: out = 16'h409D;
            12'd4058: out = 16'h4099;
            12'd4059: out = 16'h4095;
            12'd4060: out = 16'h4091;
            12'd4061: out = 16'h408D;
            12'd4062: out = 16'h4089;
            12'd4063: out = 16'h4085;
            12'd4064: out = 16'h4081;
            12'd4065: out = 16'h407D;
            12'd4066: out = 16'h4079;
            12'd4067: out = 16'h4075;
            12'd4068: out = 16'h4071;
            12'd4069: out = 16'h406D;
            12'd4070: out = 16'h4069;
            12'd4071: out = 16'h4065;
            12'd4072: out = 16'h4061;
            12'd4073: out = 16'h405D;
            12'd4074: out = 16'h4058;
            12'd4075: out = 16'h4054;
            12'd4076: out = 16'h4050;
            12'd4077: out = 16'h404C;
            12'd4078: out = 16'h4048;
            12'd4079: out = 16'h4044;
            12'd4080: out = 16'h4040;
            12'd4081: out = 16'h403C;
            12'd4082: out = 16'h4038;
            12'd4083: out = 16'h4034;
            12'd4084: out = 16'h4030;
            12'd4085: out = 16'h402C;
            12'd4086: out = 16'h4028;
            12'd4087: out = 16'h4024;
            12'd4088: out = 16'h4020;
            12'd4089: out = 16'h401C;
            12'd4090: out = 16'h4018;
            12'd4091: out = 16'h4014;
            12'd4092: out = 16'h4010;
            12'd4093: out = 16'h400C;
            12'd4094: out = 16'h4008;
            12'd4095: out = 16'h4004;
            default:  out = 16'h0000;
        endcase
    end
endmodule
