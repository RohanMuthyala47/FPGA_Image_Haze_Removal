// Atmospheric Light Estimation Module
module ALE(
    input         clk,
    input         rst,
    
    input         input_is_valid,   // Input data valid signal
    
    input [23:0]  input_pixel_1,
    input [23:0]  input_pixel_2,
    input [23:0]  input_pixel_3,
    input [23:0]  input_pixel_4,
    input [23:0]  input_pixel_5,
    input [23:0]  input_pixel_6,
    input [23:0]  input_pixel_7,
    input [23:0]  input_pixel_8,
    input [23:0]  input_pixel_9,    // 3x3 window input
    
    output [7:0]  A_R,
    output [7:0]  A_G,
    output [7:0]  A_B,              // Atmospheric Light Values
    
    output [15:0] Inv_A_R,
    output [15:0] Inv_A_G,
    output [15:0] Inv_A_B,          // Inverse Atmospheric Light Values
    
    output        output_is_valid   // Output data valid signal
);
    
    // Minimum of 9 - R/G/B channels (output wires)
    wire [7:0] minimum_red, minimum_green, minimum_blue;
    
    // Pipeline Registers (Stage 1)
    reg [7:0] minimum_red_P, minimum_green_P, minimum_blue_P;
    
    always @(posedge clk) begin
        if(rst) begin
            minimum_red_P <= 8'd0;
            minimum_green_P <= 8'd0;
            minimum_blue_P <= 8'd0;
        end
        else begin
            minimum_red_P <= minimum_red;
            minimum_green_P <= minimum_green;
            minimum_blue_P <= minimum_blue;
        end
    end
    
    wire [7:0] Dark_channel;
    
    // LUT outputs
    wire [15:0] LUT_Inv_AR, LUT_Inv_AG, LUT_Inv_AB;
    
    wire [7:0] Dark_channel_Red, Dark_channel_Green, Dark_channel_Blue;
    
    // Pipeline Registers (Stage 2)
    reg [7:0]  Dark_channel_P;
    reg [7:0]  AR_P, AG_P, AB_P;
    reg [15:0] Inv_AR_P, Inv_AG_P, Inv_AB_P;
    
    assign Dark_channel_Red = (Dark_channel > Dark_channel_P) ? (minimum_red_P * 7) >> 3 : AR_P;
    assign Dark_channel_Green = (Dark_channel > Dark_channel_P) ? (minimum_green_P * 7) >> 3 : AG_P;
    assign Dark_channel_Blue = (Dark_channel > Dark_channel_P) ? (minimum_blue_P * 7) >> 3 : AB_P;
    
    always @(posedge clk) begin
        if(rst) begin
            Dark_channel_P <= 8'd0;
            
            AR_P <= 8'd0;
            AG_P <= 8'd0;
            AB_P <= 8'd0;
            
            Inv_AR_P <= 16'd0;
            Inv_AG_P <= 16'd0;
            Inv_AB_P <= 16'd0;
        end
        else begin
            Dark_channel_P <= (Dark_channel > Dark_channel_P) ? Dark_channel : Dark_channel_P;
            
            AR_P <= Dark_channel_Red;
            AG_P <= Dark_channel_Green;
            AB_P <= Dark_channel_Blue;
            
            Inv_AR_P <= LUT_Inv_AR;
            Inv_AG_P <= LUT_Inv_AG;
            Inv_AB_P <= LUT_Inv_AB;
        end
    end
    
    // Delay the valid signal by 2 clock cycles
    reg Stage_1_valid, Stage_2_valid;
    always @(posedge clk)
    begin
        if(rst) begin
            Stage_1_valid <= 0;
            Stage_2_valid <= 0;
        end
        else begin
            Stage_1_valid <= input_is_valid;
            Stage_2_valid <= Stage_1_valid;
        end
    end
    
    // Output wire assignments
    assign A_R = AR_P;
    assign A_G = AG_P;
    assign A_B = AB_P;
    
    assign Inv_A_R = Inv_AR_P;
    assign Inv_A_G = Inv_AG_P;
    assign Inv_A_B = Inv_AB_P;
    
    assign output_is_valid = Stage_2_valid;

/////////////////////////////////////////////////////////////////////////////////
// BLOCK DECLARATIONS
/////////////////////////////////////////////////////////////////////////////////

    // Find the minimum of each color channel inputs
    ALE_Minimum_9 Red (
        .input_pixel_1(input_pixel_1[23:16]),
        .input_pixel_2(input_pixel_2[23:16]),
        .input_pixel_3(input_pixel_3[23:16]),
        .input_pixel_4(input_pixel_4[23:16]),
        .input_pixel_5(input_pixel_5[23:16]),
        .input_pixel_6(input_pixel_6[23:16]),
        .input_pixel_7(input_pixel_7[23:16]),
        .input_pixel_8(input_pixel_8[23:16]),
        .input_pixel_9(input_pixel_9[23:16]),
        .minimum_pixel(minimum_red)
    );
    
    ALE_Minimum_9 Green (
        .input_pixel_1(input_pixel_1[15:8]),
        .input_pixel_2(input_pixel_2[15:8]),
        .input_pixel_3(input_pixel_3[15:8]),
        .input_pixel_4(input_pixel_4[15:8]),
        .input_pixel_5(input_pixel_5[15:8]),
        .input_pixel_6(input_pixel_6[15:8]),
        .input_pixel_7(input_pixel_7[15:8]),
        .input_pixel_8(input_pixel_8[15:8]),
        .input_pixel_9(input_pixel_9[15:8]),
        .minimum_pixel(minimum_green)
    );
    
    ALE_Minimum_9 Blue (
        .input_pixel_1(input_pixel_1[7:0]),
        .input_pixel_2(input_pixel_2[7:0]),
        .input_pixel_3(input_pixel_3[7:0]),
        .input_pixel_4(input_pixel_4[7:0]),
        .input_pixel_5(input_pixel_5[7:0]),
        .input_pixel_6(input_pixel_6[7:0]),
        .input_pixel_7(input_pixel_7[7:0]),
        .input_pixel_8(input_pixel_8[7:0]),
        .input_pixel_9(input_pixel_9[7:0]),
        .minimum_pixel(minimum_blue)
    );
    
    // Calculate minimum among the three channels to get dark channel
    ALE_Minimum_3 Dark_Channel(
        .a(minimum_red_P), .b(minimum_green_P), .c(minimum_blue_P),
        .minimum(Dark_channel)
    );
    
    // Look-Up Tables to output the reciprocal of the atmospheric light value in Q0.16 format
    ATM_LUT Inverse_Red(
        .in_val(Dark_channel_Red),
        .out_val(LUT_Inv_AR)
    );
    
    ATM_LUT Inverse_Green(
        .in_val(Dark_channel_Green),
        .out_val(LUT_Inv_AG)
    );
    
    ATM_LUT Inverse_Blue(
        .in_val(Dark_channel_Blue),
        .out_val(LUT_Inv_AB)
    );
    
endmodule
