module Transmission_Reciprocal_LUT (
    input  [7:0] in,      // Q0.8 input (unsigned Q0.8 value ranging from 0 to 0.65)
    output reg [7:0] out  // Q2.6 reciprocal output (unsigned, 8-bit)
);

    always @(*) begin
        case(in)
            8'd  0: out = 8'h40;
            8'd  1: out = 8'h40;
            8'd  2: out = 8'h41;
            8'd  3: out = 8'h41;
            8'd  4: out = 8'h41;
            8'd  5: out = 8'h41;
            8'd  6: out = 8'h42;
            8'd  7: out = 8'h42;
            8'd  8: out = 8'h42;
            8'd  9: out = 8'h42;
            8'd 10: out = 8'h43;
            8'd 11: out = 8'h43;
            8'd 12: out = 8'h43;
            8'd 13: out = 8'h43;
            8'd 14: out = 8'h44;
            8'd 15: out = 8'h44;
            8'd 16: out = 8'h44;
            8'd 17: out = 8'h45;
            8'd 18: out = 8'h45;
            8'd 19: out = 8'h45;
            8'd 20: out = 8'h45;
            8'd 21: out = 8'h46;
            8'd 22: out = 8'h46;
            8'd 23: out = 8'h46;
            8'd 24: out = 8'h47;
            8'd 25: out = 8'h47;
            8'd 26: out = 8'h47;
            8'd 27: out = 8'h48;
            8'd 28: out = 8'h48;
            8'd 29: out = 8'h48;
            8'd 30: out = 8'h48;
            8'd 31: out = 8'h49;
            8'd 32: out = 8'h49;
            8'd 33: out = 8'h49;
            8'd 34: out = 8'h4A;
            8'd 35: out = 8'h4A;
            8'd 36: out = 8'h4A;
            8'd 37: out = 8'h4B;
            8'd 38: out = 8'h4B;
            8'd 39: out = 8'h4C;
            8'd 40: out = 8'h4C;
            8'd 41: out = 8'h4C;
            8'd 42: out = 8'h4D;
            8'd 43: out = 8'h4D;
            8'd 44: out = 8'h4D;
            8'd 45: out = 8'h4E;
            8'd 46: out = 8'h4E;
            8'd 47: out = 8'h4E;
            8'd 48: out = 8'h4F;
            8'd 49: out = 8'h4F;
            8'd 50: out = 8'h50;
            8'd 51: out = 8'h50;
            8'd 52: out = 8'h50;
            8'd 53: out = 8'h51;
            8'd 54: out = 8'h51;
            8'd 55: out = 8'h52;
            8'd 56: out = 8'h52;
            8'd 57: out = 8'h52;
            8'd 58: out = 8'h53;
            8'd 59: out = 8'h53;
            8'd 60: out = 8'h54;
            8'd 61: out = 8'h54;
            8'd 62: out = 8'h54;
            8'd 63: out = 8'h55;
            8'd 64: out = 8'h55;
            8'd 65: out = 8'h56;
            8'd 66: out = 8'h56;
            8'd 67: out = 8'h57;
            8'd 68: out = 8'h57;
            8'd 69: out = 8'h58;
            8'd 70: out = 8'h58;
            8'd 71: out = 8'h59;
            8'd 72: out = 8'h59;
            8'd 73: out = 8'h5A;
            8'd 74: out = 8'h5A;
            8'd 75: out = 8'h5B;
            8'd 76: out = 8'h5B;
            8'd 77: out = 8'h5C;
            8'd 78: out = 8'h5C;
            8'd 79: out = 8'h5D;
            8'd 80: out = 8'h5D;
            8'd 81: out = 8'h5E;
            8'd 82: out = 8'h5E;
            8'd 83: out = 8'h5F;
            8'd 84: out = 8'h5F;
            8'd 85: out = 8'h60;
            8'd 86: out = 8'h60;
            8'd 87: out = 8'h61;
            8'd 88: out = 8'h62;
            8'd 89: out = 8'h62;
            8'd 90: out = 8'h63;
            8'd 91: out = 8'h63;
            8'd 92: out = 8'h64;
            8'd 93: out = 8'h65;
            8'd 94: out = 8'h65;
            8'd 95: out = 8'h66;
            8'd 96: out = 8'h66;
            8'd 97: out = 8'h67;
            8'd 98: out = 8'h68;
            8'd 99: out = 8'h68;
            8'd100: out = 8'h69;
            8'd101: out = 8'h6A;
            8'd102: out = 8'h6A;
            8'd103: out = 8'h6B;
            8'd104: out = 8'h6C;
            8'd105: out = 8'h6D;
            8'd106: out = 8'h6D;
            8'd107: out = 8'h6E;
            8'd108: out = 8'h6F;
            8'd109: out = 8'h6F;
            8'd110: out = 8'h70;
            8'd111: out = 8'h71;
            8'd112: out = 8'h72;
            8'd113: out = 8'h73;
            8'd114: out = 8'h73;
            8'd115: out = 8'h74;
            8'd116: out = 8'h75;
            8'd117: out = 8'h76;
            8'd118: out = 8'h77;
            8'd119: out = 8'h78;
            8'd120: out = 8'h78;
            8'd121: out = 8'h79;
            8'd122: out = 8'h7A;
            8'd123: out = 8'h7B;
            8'd124: out = 8'h7C;
            8'd125: out = 8'h7D;
            8'd126: out = 8'h7E;
            8'd127: out = 8'h7F;
            8'd128: out = 8'h80;
            8'd129: out = 8'h81;
            8'd130: out = 8'h82;
            8'd131: out = 8'h83;
            8'd132: out = 8'h84;
            8'd133: out = 8'h85;
            8'd134: out = 8'h86;
            8'd135: out = 8'h87;
            8'd136: out = 8'h89;
            8'd137: out = 8'h8A;
            8'd138: out = 8'h8B;
            8'd139: out = 8'h8C;
            8'd140: out = 8'h8D;
            8'd141: out = 8'h8E;
            8'd142: out = 8'h90;
            8'd143: out = 8'h91;
            8'd144: out = 8'h92;
            8'd145: out = 8'h94;
            8'd146: out = 8'h95;
            8'd147: out = 8'h96;
            8'd148: out = 8'h98;
            8'd149: out = 8'h99;
            8'd150: out = 8'h9B;
            8'd151: out = 8'h9C;
            8'd152: out = 8'h9E;
            8'd153: out = 8'h9F;
            8'd154: out = 8'hA1;
            8'd155: out = 8'hA2;
            8'd156: out = 8'hA4;
            8'd157: out = 8'hA5;
            8'd158: out = 8'hA7;
            8'd159: out = 8'hA9;
            8'd160: out = 8'hAB;
            8'd161: out = 8'hAC;
            8'd162: out = 8'hAE;
            8'd163: out = 8'hB0;
            8'd164: out = 8'hB2;
            8'd165: out = 8'hB4;
            8'd166: out = 8'hB6;
            default: out = 8'hB8;
        endcase
    end
endmodule
