// Look Up Tables for applying saturation correction

module LUT_03 (
    input       [7:0] x,
    output reg [15:0] y // Q3.13 format
);

    always @(*) begin
        case (x)
            8'd0  : y = 16'd0;  // 0^0.3 ~= 0.000000
            8'd1  : y = 16'd8192;  // 1^0.3 ~= 1.000000
            8'd2  : y = 16'd10086;  // 2^0.3 ~= 1.231144
            8'd3  : y = 16'd11390;  // 3^0.3 ~= 1.390389
            8'd4  : y = 16'd12417;  // 4^0.3 ~= 1.515717
            8'd5  : y = 16'd13276;  // 5^0.3 ~= 1.620657
            8'd6  : y = 16'd14023;  // 6^0.3 ~= 1.711770
            8'd7  : y = 16'd14687;  // 7^0.3 ~= 1.792790
            8'd8  : y = 16'd15287;  // 8^0.3 ~= 1.866066
            8'd9  : y = 16'd15837;  // 9^0.3 ~= 1.933182
            8'd10 : y = 16'd16345;  // 10^0.3 ~= 1.995262
            8'd11 : y = 16'd16819;  // 11^0.3 ~= 2.053136
            8'd12 : y = 16'd17264;  // 12^0.3 ~= 2.107436
            8'd13 : y = 16'd17684;  // 13^0.3 ~= 2.158654
            8'd14 : y = 16'd18081;  // 14^0.3 ~= 2.207183
            8'd15 : y = 16'd18459;  // 15^0.3 ~= 2.253343
            8'd16 : y = 16'd18820;  // 16^0.3 ~= 2.297397
            8'd17 : y = 16'd19166;  // 17^0.3 ~= 2.339563
            8'd18 : y = 16'd19497;  // 18^0.3 ~= 2.380026
            8'd19 : y = 16'd19816;  // 19^0.3 ~= 2.418945
            8'd20 : y = 16'd20123;  // 20^0.3 ~= 2.456456
            8'd21 : y = 16'd20420;  // 21^0.3 ~= 2.492676
            8'd22 : y = 16'd20707;  // 22^0.3 ~= 2.527707
            8'd23 : y = 16'd20985;  // 23^0.3 ~= 2.561642
            8'd24 : y = 16'd21255;  // 24^0.3 ~= 2.594558
            8'd25 : y = 16'd21517;  // 25^0.3 ~= 2.626528
            8'd26 : y = 16'd21771;  // 26^0.3 ~= 2.657615
            8'd27 : y = 16'd22019;  // 27^0.3 ~= 2.687875
            8'd28 : y = 16'd22261;  // 28^0.3 ~= 2.717361
            8'd29 : y = 16'd22496;  // 29^0.3 ~= 2.746119
            8'd30 : y = 16'd22726;  // 30^0.3 ~= 2.774191
            8'd31 : y = 16'd22951;  // 31^0.3 ~= 2.801615
            8'd32 : y = 16'd23170;  // 32^0.3 ~= 2.828427
            8'd33 : y = 16'd23385;  // 33^0.3 ~= 2.854659
            8'd34 : y = 16'd23596;  // 34^0.3 ~= 2.880339
            8'd35 : y = 16'd23802;  // 35^0.3 ~= 2.905497
            8'd36 : y = 16'd24004;  // 36^0.3 ~= 2.930156
            8'd37 : y = 16'd24202;  // 37^0.3 ~= 2.954340
            8'd38 : y = 16'd24396;  // 38^0.3 ~= 2.978071
            8'd39 : y = 16'd24587;  // 39^0.3 ~= 3.001369
            8'd40 : y = 16'd24775;  // 40^0.3 ~= 3.024252
            8'd41 : y = 16'd24959;  // 41^0.3 ~= 3.046738
            8'd42 : y = 16'd25140;  // 42^0.3 ~= 3.068844
            8'd43 : y = 16'd25318;  // 43^0.3 ~= 3.090584
            8'd44 : y = 16'd25493;  // 44^0.3 ~= 3.111973
            8'd45 : y = 16'd25666;  // 45^0.3 ~= 3.133024
            8'd46 : y = 16'd25836;  // 46^0.3 ~= 3.153751
            8'd47 : y = 16'd26003;  // 47^0.3 ~= 3.174164
            8'd48 : y = 16'd26168;  // 48^0.3 ~= 3.194276
            8'd49 : y = 16'd26330;  // 49^0.3 ~= 3.214096
            8'd50 : y = 16'd26490;  // 50^0.3 ~= 3.233635
            8'd51 : y = 16'd26648;  // 51^0.3 ~= 3.252903
            8'd52 : y = 16'd26803;  // 52^0.3 ~= 3.271907
            8'd53 : y = 16'd26957;  // 53^0.3 ~= 3.290658
            8'd54 : y = 16'd27109;  // 54^0.3 ~= 3.309163
            8'd55 : y = 16'd27258;  // 55^0.3 ~= 3.327429
            8'd56 : y = 16'd27406;  // 56^0.3 ~= 3.345464
            8'd57 : y = 16'd27552;  // 57^0.3 ~= 3.363276
            8'd58 : y = 16'd27696;  // 58^0.3 ~= 3.380869
            8'd59 : y = 16'd27838;  // 59^0.3 ~= 3.398252
            8'd60 : y = 16'd27979;  // 60^0.3 ~= 3.415430
            8'd61 : y = 16'd28118;  // 61^0.3 ~= 3.432408
            8'd62 : y = 16'd28256;  // 62^0.3 ~= 3.449193
            8'd63 : y = 16'd28392;  // 63^0.3 ~= 3.465789
            8'd64 : y = 16'd28526;  // 64^0.3 ~= 3.482202
            8'd65 : y = 16'd28659;  // 65^0.3 ~= 3.498437
            8'd66 : y = 16'd28791;  // 66^0.3 ~= 3.514497
            8'd67 : y = 16'd28921;  // 67^0.3 ~= 3.530388
            8'd68 : y = 16'd29050;  // 68^0.3 ~= 3.546114
            8'd69 : y = 16'd29177;  // 69^0.3 ~= 3.561679
            8'd70 : y = 16'd29303;  // 70^0.3 ~= 3.577086
            8'd71 : y = 16'd29428;  // 71^0.3 ~= 3.592341
            8'd72 : y = 16'd29552;  // 72^0.3 ~= 3.607445
            8'd73 : y = 16'd29675;  // 73^0.3 ~= 3.622404
            8'd74 : y = 16'd29796;  // 74^0.3 ~= 3.637220
            8'd75 : y = 16'd29916;  // 75^0.3 ~= 3.651896
            8'd76 : y = 16'd30035;  // 76^0.3 ~= 3.666436
            8'd77 : y = 16'd30153;  // 77^0.3 ~= 3.680842
            8'd78 : y = 16'd30270;  // 78^0.3 ~= 3.695119
            8'd79 : y = 16'd30386;  // 79^0.3 ~= 3.709267
            8'd80 : y = 16'd30501;  // 80^0.3 ~= 3.723291
            8'd81 : y = 16'd30615;  // 81^0.3 ~= 3.737193
            8'd82 : y = 16'd30728;  // 82^0.3 ~= 3.750975
            8'd83 : y = 16'd30840;  // 83^0.3 ~= 3.764640
            8'd84 : y = 16'd30951;  // 84^0.3 ~= 3.778190
            8'd85 : y = 16'd31061;  // 85^0.3 ~= 3.791628
            8'd86 : y = 16'd31170;  // 86^0.3 ~= 3.804955
            8'd87 : y = 16'd31278;  // 87^0.3 ~= 3.818175
            8'd88 : y = 16'd31386;  // 88^0.3 ~= 3.831288
            8'd89 : y = 16'd31492;  // 89^0.3 ~= 3.844298
            8'd90 : y = 16'd31598;  // 90^0.3 ~= 3.857205
            8'd91 : y = 16'd31703;  // 91^0.3 ~= 3.870013
            8'd92 : y = 16'd31807;  // 92^0.3 ~= 3.882722
            8'd93 : y = 16'd31911;  // 93^0.3 ~= 3.895336
            8'd94 : y = 16'd32013;  // 94^0.3 ~= 3.907854
            8'd95 : y = 16'd32115;  // 95^0.3 ~= 3.920280
            8'd96 : y = 16'd32216;  // 96^0.3 ~= 3.932614
            8'd97 : y = 16'd32316;  // 97^0.3 ~= 3.944859
            8'd98 : y = 16'd32416;  // 98^0.3 ~= 3.957016
            8'd99 : y = 16'd32515;  // 99^0.3 ~= 3.969086
            8'd100: y = 16'd32613;  // 100^0.3 ~= 3.981072
            8'd101: y = 16'd32710;  // 101^0.3 ~= 3.992973
            8'd102: y = 16'd32807;  // 102^0.3 ~= 4.004793
            8'd103: y = 16'd32903;  // 103^0.3 ~= 4.016531
            8'd104: y = 16'd32999;  // 104^0.3 ~= 4.028191
            8'd105: y = 16'd33094;  // 105^0.3 ~= 4.039771
            8'd106: y = 16'd33188;  // 106^0.3 ~= 4.051275
            8'd107: y = 16'd33282;  // 107^0.3 ~= 4.062704
            8'd108: y = 16'd33375;  // 108^0.3 ~= 4.074057
            8'd109: y = 16'd33467;  // 109^0.3 ~= 4.085338
            8'd110: y = 16'd33559;  // 110^0.3 ~= 4.096546
            8'd111: y = 16'd33650;  // 111^0.3 ~= 4.107683
            8'd112: y = 16'd33741;  // 112^0.3 ~= 4.118750
            8'd113: y = 16'd33831;  // 113^0.3 ~= 4.129748
            8'd114: y = 16'd33920;  // 114^0.3 ~= 4.140678
            8'd115: y = 16'd34009;  // 115^0.3 ~= 4.151541
            8'd116: y = 16'd34098;  // 116^0.3 ~= 4.162339
            8'd117: y = 16'd34186;  // 117^0.3 ~= 4.173071
            8'd118: y = 16'd34273;  // 118^0.3 ~= 4.183739
            8'd119: y = 16'd34360;  // 119^0.3 ~= 4.194344
            8'd120: y = 16'd34446;  // 120^0.3 ~= 4.204887
            8'd121: y = 16'd34532;  // 121^0.3 ~= 4.215369
            8'd122: y = 16'd34618;  // 122^0.3 ~= 4.225790
            8'd123: y = 16'd34703;  // 123^0.3 ~= 4.236152
            8'd124: y = 16'd34787;  // 124^0.3 ~= 4.246455
            8'd125: y = 16'd34871;  // 125^0.3 ~= 4.256700
            8'd126: y = 16'd34954;  // 126^0.3 ~= 4.266887
            8'd127: y = 16'd35037;  // 127^0.3 ~= 4.277018
            8'd128: y = 16'd35120;  // 128^0.3 ~= 4.287094
            8'd129: y = 16'd35202;  // 129^0.3 ~= 4.297114
            8'd130: y = 16'd35284;  // 130^0.3 ~= 4.307081
            8'd131: y = 16'd35365;  // 131^0.3 ~= 4.316993
            8'd132: y = 16'd35446;  // 132^0.3 ~= 4.326853
            8'd133: y = 16'd35526;  // 133^0.3 ~= 4.336661
            8'd134: y = 16'd35606;  // 134^0.3 ~= 4.346417
            8'd135: y = 16'd35685;  // 135^0.3 ~= 4.356123
            8'd136: y = 16'd35764;  // 136^0.3 ~= 4.365778
            8'd137: y = 16'd35843;  // 137^0.3 ~= 4.375384
            8'd138: y = 16'd35921;  // 138^0.3 ~= 4.384941
            8'd139: y = 16'd35999;  // 139^0.3 ~= 4.394449
            8'd140: y = 16'd36077;  // 140^0.3 ~= 4.403910
            8'd141: y = 16'd36154;  // 141^0.3 ~= 4.413323
            8'd142: y = 16'd36231;  // 142^0.3 ~= 4.422690
            8'd143: y = 16'd36307;  // 143^0.3 ~= 4.432011
            8'd144: y = 16'd36383;  // 144^0.3 ~= 4.441286
            8'd145: y = 16'd36459;  // 145^0.3 ~= 4.450516
            8'd146: y = 16'd36534;  // 146^0.3 ~= 4.459702
            8'd147: y = 16'd36609;  // 147^0.3 ~= 4.468844
            8'd148: y = 16'd36683;  // 148^0.3 ~= 4.477943
            8'd149: y = 16'd36757;  // 149^0.3 ~= 4.486998
            8'd150: y = 16'd36831;  // 150^0.3 ~= 4.496011
            8'd151: y = 16'd36905;  // 151^0.3 ~= 4.504982
            8'd152: y = 16'd36978;  // 152^0.3 ~= 4.513912
            8'd153: y = 16'd37051;  // 153^0.3 ~= 4.522800
            8'd154: y = 16'd37123;  // 154^0.3 ~= 4.531649
            8'd155: y = 16'd37195;  // 155^0.3 ~= 4.540456
            8'd156: y = 16'd37267;  // 156^0.3 ~= 4.549225
            8'd157: y = 16'd37339;  // 157^0.3 ~= 4.557954
            8'd158: y = 16'd37410;  // 158^0.3 ~= 4.566644
            8'd159: y = 16'd37481;  // 159^0.3 ~= 4.575295
            8'd160: y = 16'd37551;  // 160^0.3 ~= 4.583909
            8'd161: y = 16'd37622;  // 161^0.3 ~= 4.592485
            8'd162: y = 16'd37692;  // 162^0.3 ~= 4.601024
            8'd163: y = 16'd37761;  // 163^0.3 ~= 4.609526
            8'd164: y = 16'd37831;  // 164^0.3 ~= 4.617992
            8'd165: y = 16'd37900;  // 165^0.3 ~= 4.626421
            8'd166: y = 16'd37968;  // 166^0.3 ~= 4.634815
            8'd167: y = 16'd38037;  // 167^0.3 ~= 4.643174
            8'd168: y = 16'd38105;  // 168^0.3 ~= 4.651497
            8'd169: y = 16'd38173;  // 169^0.3 ~= 4.659786
            8'd170: y = 16'd38241;  // 170^0.3 ~= 4.668041
            8'd171: y = 16'd38308;  // 171^0.3 ~= 4.676262
            8'd172: y = 16'd38375;  // 172^0.3 ~= 4.684449
            8'd173: y = 16'd38442;  // 173^0.3 ~= 4.692603
            8'd174: y = 16'd38508;  // 174^0.3 ~= 4.700724
            8'd175: y = 16'd38575;  // 175^0.3 ~= 4.708813
            8'd176: y = 16'd38641;  // 176^0.3 ~= 4.716869
            8'd177: y = 16'd38706;  // 177^0.3 ~= 4.724893
            8'd178: y = 16'd38772;  // 178^0.3 ~= 4.732886
            8'd179: y = 16'd38837;  // 179^0.3 ~= 4.740847
            8'd180: y = 16'd38902;  // 180^0.3 ~= 4.748777
            8'd181: y = 16'd38967;  // 181^0.3 ~= 4.756676
            8'd182: y = 16'd39031;  // 182^0.3 ~= 4.764545
            8'd183: y = 16'd39095;  // 183^0.3 ~= 4.772383
            8'd184: y = 16'd39159;  // 184^0.3 ~= 4.780192
            8'd185: y = 16'd39223;  // 185^0.3 ~= 4.787971
            8'd186: y = 16'd39287;  // 186^0.3 ~= 4.795721
            8'd187: y = 16'd39350;  // 187^0.3 ~= 4.803441
            8'd188: y = 16'd39413;  // 188^0.3 ~= 4.811133
            8'd189: y = 16'd39476;  // 189^0.3 ~= 4.818796
            8'd190: y = 16'd39538;  // 190^0.3 ~= 4.826431
            8'd191: y = 16'd39600;  // 191^0.3 ~= 4.834037
            8'd192: y = 16'd39663;  // 192^0.3 ~= 4.841616
            8'd193: y = 16'd39724;  // 193^0.3 ~= 4.849168
            8'd194: y = 16'd39786;  // 194^0.3 ~= 4.856692
            8'd195: y = 16'd39847;  // 195^0.3 ~= 4.864188
            8'd196: y = 16'd39909;  // 196^0.3 ~= 4.871658
            8'd197: y = 16'd39970;  // 197^0.3 ~= 4.879102
            8'd198: y = 16'd40030;  // 198^0.3 ~= 4.886519
            8'd199: y = 16'd40091;  // 199^0.3 ~= 4.893909
            8'd200: y = 16'd40151;  // 200^0.3 ~= 4.901274
            8'd201: y = 16'd40211;  // 201^0.3 ~= 4.908613
            8'd202: y = 16'd40271;  // 202^0.3 ~= 4.915927
            8'd203: y = 16'd40331;  // 203^0.3 ~= 4.923215
            8'd204: y = 16'd40390;  // 204^0.3 ~= 4.930478
            8'd205: y = 16'd40450;  // 205^0.3 ~= 4.937717
            8'd206: y = 16'd40509;  // 206^0.3 ~= 4.944930
            8'd207: y = 16'd40568;  // 207^0.3 ~= 4.952119
            8'd208: y = 16'd40626;  // 208^0.3 ~= 4.959284
            8'd209: y = 16'd40685;  // 209^0.3 ~= 4.966425
            8'd210: y = 16'd40743;  // 210^0.3 ~= 4.973542
            8'd211: y = 16'd40801;  // 211^0.3 ~= 4.980635
            8'd212: y = 16'd40859;  // 212^0.3 ~= 4.987705
            8'd213: y = 16'd40917;  // 213^0.3 ~= 4.994751
            8'd214: y = 16'd40975;  // 214^0.3 ~= 5.001775
            8'd215: y = 16'd41032;  // 215^0.3 ~= 5.008775
            8'd216: y = 16'd41089;  // 216^0.3 ~= 5.015753
            8'd217: y = 16'd41146;  // 217^0.3 ~= 5.022708
            8'd218: y = 16'd41203;  // 218^0.3 ~= 5.029641
            8'd219: y = 16'd41259;  // 219^0.3 ~= 5.036551
            8'd220: y = 16'd41316;  // 220^0.3 ~= 5.043439
            8'd221: y = 16'd41372;  // 221^0.3 ~= 5.050306
            8'd222: y = 16'd41428;  // 222^0.3 ~= 5.057151
            8'd223: y = 16'd41484;  // 223^0.3 ~= 5.063974
            8'd224: y = 16'd41540;  // 224^0.3 ~= 5.070776
            8'd225: y = 16'd41595;  // 225^0.3 ~= 5.077556
            8'd226: y = 16'd41651;  // 226^0.3 ~= 5.084316
            8'd227: y = 16'd41706;  // 227^0.3 ~= 5.091055
            8'd228: y = 16'd41761;  // 228^0.3 ~= 5.097773
            8'd229: y = 16'd41816;  // 229^0.3 ~= 5.104470
            8'd230: y = 16'd41871;  // 230^0.3 ~= 5.111147
            8'd231: y = 16'd41925;  // 231^0.3 ~= 5.117803
            8'd232: y = 16'd41979;  // 232^0.3 ~= 5.124440
            8'd233: y = 16'd42034;  // 233^0.3 ~= 5.131056
            8'd234: y = 16'd42088;  // 234^0.3 ~= 5.137653
            8'd235: y = 16'd42142;  // 235^0.3 ~= 5.144230
            8'd236: y = 16'd42195;  // 236^0.3 ~= 5.150787
            8'd237: y = 16'd42249;  // 237^0.3 ~= 5.157325
            8'd238: y = 16'd42302;  // 238^0.3 ~= 5.163844
            8'd239: y = 16'd42355;  // 239^0.3 ~= 5.170343
            8'd240: y = 16'd42409;  // 240^0.3 ~= 5.176824
            8'd241: y = 16'd42461;  // 241^0.3 ~= 5.183285
            8'd242: y = 16'd42514;  // 242^0.3 ~= 5.189728
            8'd243: y = 16'd42567;  // 243^0.3 ~= 5.196152
            8'd244: y = 16'd42619;  // 244^0.3 ~= 5.202558
            8'd245: y = 16'd42672;  // 245^0.3 ~= 5.208946
            8'd246: y = 16'd42724;  // 246^0.3 ~= 5.215315
            8'd247: y = 16'd42776;  // 247^0.3 ~= 5.221666
            8'd248: y = 16'd42828;  // 248^0.3 ~= 5.227999
            8'd249: y = 16'd42880;  // 249^0.3 ~= 5.234314
            8'd250: y = 16'd42931;  // 250^0.3 ~= 5.240612
            8'd251: y = 16'd42983;  // 251^0.3 ~= 5.246892
            8'd252: y = 16'd43034;  // 252^0.3 ~= 5.253154
            8'd253: y = 16'd43085;  // 253^0.3 ~= 5.259399
            8'd254: y = 16'd43136;  // 254^0.3 ~= 5.265627
            8'd255: y = 16'd43187;  // 255^0.3 ~= 5.271838
            default: y = 16'd0;
        endcase
    end
endmodule

module LUT_07 (
    input       [7:0] x,
    output reg [15:0] y // Q6.10 format
);

    always @(*) begin
        case (x)
            8'd0  : y = 16'd0;  // 0^0.7 ~= 0.000000
            8'd1  : y = 16'd1024;  // 1^0.7 ~= 1.000000
            8'd2  : y = 16'd1663;  // 2^0.7 ~= 1.624505
            8'd3  : y = 16'd2209;  // 3^0.7 ~= 2.157669
            8'd4  : y = 16'd2702;  // 4^0.7 ~= 2.639016
            8'd5  : y = 16'd3159;  // 5^0.7 ~= 3.085169
            8'd6  : y = 16'd3589;  // 6^0.7 ~= 3.505144
            8'd7  : y = 16'd3998;  // 7^0.7 ~= 3.904529
            8'd8  : y = 16'd4390;  // 8^0.7 ~= 4.287094
            8'd9  : y = 16'd4767;  // 9^0.7 ~= 4.655537
            8'd10 : y = 16'd5132;  // 10^0.7 ~= 5.011872
            8'd11 : y = 16'd5486;  // 11^0.7 ~= 5.357657
            8'd12 : y = 16'd5831;  // 12^0.7 ~= 5.694123
            8'd13 : y = 16'd6167;  // 13^0.7 ~= 6.022272
            8'd14 : y = 16'd6495;  // 14^0.7 ~= 6.342926
            8'd15 : y = 16'd6817;  // 15^0.7 ~= 6.656775
            8'd16 : y = 16'd7132;  // 16^0.7 ~= 6.964405
            8'd17 : y = 16'd7441;  // 17^0.7 ~= 7.266315
            8'd18 : y = 16'd7744;  // 18^0.7 ~= 7.562942
            8'd19 : y = 16'd8043;  // 19^0.7 ~= 7.854662
            8'd20 : y = 16'd8337;  // 20^0.7 ~= 8.141811
            8'd21 : y = 16'd8627;  // 21^0.7 ~= 8.424682
            8'd22 : y = 16'd8912;  // 22^0.7 ~= 8.703539
            8'd23 : y = 16'd9194;  // 23^0.7 ~= 8.978618
            8'd24 : y = 16'd9472;  // 24^0.7 ~= 9.250131
            8'd25 : y = 16'd9747;  // 25^0.7 ~= 9.518270
            8'd26 : y = 16'd10018;  // 26^0.7 ~= 9.783209
            8'd27 : y = 16'd10286;  // 27^0.7 ~= 10.045109
            8'd28 : y = 16'd10551;  // 28^0.7 ~= 10.304113
            8'd29 : y = 16'd10814;  // 29^0.7 ~= 10.560357
            8'd30 : y = 16'd11073;  // 30^0.7 ~= 10.813963
            8'd31 : y = 16'd11331;  // 31^0.7 ~= 11.065045
            8'd32 : y = 16'd11585;  // 32^0.7 ~= 11.313708
            8'd33 : y = 16'd11837;  // 33^0.7 ~= 11.560051
            8'd34 : y = 16'd12087;  // 34^0.7 ~= 11.804164
            8'd35 : y = 16'd12335;  // 35^0.7 ~= 12.046132
            8'd36 : y = 16'd12581;  // 36^0.7 ~= 12.286035
            8'd37 : y = 16'd12825;  // 37^0.7 ~= 12.523947
            8'd38 : y = 16'd13066;  // 38^0.7 ~= 12.759937
            8'd39 : y = 16'd13306;  // 39^0.7 ~= 12.994071
            8'd40 : y = 16'd13544;  // 40^0.7 ~= 13.226410
            8'd41 : y = 16'd13780;  // 41^0.7 ~= 13.457014
            8'd42 : y = 16'd14014;  // 42^0.7 ~= 13.685936
            8'd43 : y = 16'd14247;  // 43^0.7 ~= 13.913229
            8'd44 : y = 16'd14478;  // 44^0.7 ~= 14.138941
            8'd45 : y = 16'd14708;  // 45^0.7 ~= 14.363119
            8'd46 : y = 16'd14936;  // 46^0.7 ~= 14.585808
            8'd47 : y = 16'd15162;  // 47^0.7 ~= 14.807049
            8'd48 : y = 16'd15388;  // 48^0.7 ~= 15.026882
            8'd49 : y = 16'd15611;  // 49^0.7 ~= 15.245345
            8'd50 : y = 16'd15834;  // 50^0.7 ~= 15.462475
            8'd51 : y = 16'd16055;  // 51^0.7 ~= 15.678306
            8'd52 : y = 16'd16274;  // 52^0.7 ~= 15.892870
            8'd53 : y = 16'd16493;  // 53^0.7 ~= 16.106201
            8'd54 : y = 16'd16710;  // 54^0.7 ~= 16.318327
            8'd55 : y = 16'd16926;  // 55^0.7 ~= 16.529278
            8'd56 : y = 16'd17141;  // 56^0.7 ~= 16.739081
            8'd57 : y = 16'd17355;  // 57^0.7 ~= 16.947764
            8'd58 : y = 16'd17567;  // 58^0.7 ~= 17.155350
            8'd59 : y = 16'd17779;  // 59^0.7 ~= 17.361866
            8'd60 : y = 16'd17989;  // 60^0.7 ~= 17.567335
            8'd61 : y = 16'd18198;  // 61^0.7 ~= 17.771778
            8'd62 : y = 16'd18407;  // 62^0.7 ~= 17.975219
            8'd63 : y = 16'd18614;  // 63^0.7 ~= 18.177677
            8'd64 : y = 16'd18820;  // 64^0.7 ~= 18.379174
            8'd65 : y = 16'd19026;  // 65^0.7 ~= 18.579728
            8'd66 : y = 16'd19230;  // 66^0.7 ~= 18.779359
            8'd67 : y = 16'd19434;  // 67^0.7 ~= 18.978084
            8'd68 : y = 16'd19636;  // 68^0.7 ~= 19.175921
            8'd69 : y = 16'd19838;  // 69^0.7 ~= 19.372888
            8'd70 : y = 16'd20039;  // 70^0.7 ~= 19.569000
            8'd71 : y = 16'd20239;  // 71^0.7 ~= 19.764273
            8'd72 : y = 16'd20438;  // 72^0.7 ~= 19.958723
            8'd73 : y = 16'd20636;  // 73^0.7 ~= 20.152364
            8'd74 : y = 16'd20833;  // 74^0.7 ~= 20.345211
            8'd75 : y = 16'd21030;  // 75^0.7 ~= 20.537278
            8'd76 : y = 16'd21226;  // 76^0.7 ~= 20.728578
            8'd77 : y = 16'd21421;  // 77^0.7 ~= 20.919125
            8'd78 : y = 16'd21616;  // 78^0.7 ~= 21.108930
            8'd79 : y = 16'd21809;  // 79^0.7 ~= 21.298007
            8'd80 : y = 16'd22002;  // 80^0.7 ~= 21.486367
            8'd81 : y = 16'd22194;  // 81^0.7 ~= 21.674022
            8'd82 : y = 16'd22386;  // 82^0.7 ~= 21.860984
            8'd83 : y = 16'd22576;  // 83^0.7 ~= 22.047262
            8'd84 : y = 16'd22766;  // 84^0.7 ~= 22.232869
            8'd85 : y = 16'd22956;  // 85^0.7 ~= 22.417813
            8'd86 : y = 16'd23145;  // 86^0.7 ~= 22.602106
            8'd87 : y = 16'd23333;  // 87^0.7 ~= 22.785758
            8'd88 : y = 16'd23520;  // 88^0.7 ~= 22.968777
            8'd89 : y = 16'd23707;  // 89^0.7 ~= 23.151173
            8'd90 : y = 16'd23893;  // 90^0.7 ~= 23.332956
            8'd91 : y = 16'd24078;  // 91^0.7 ~= 23.514133
            8'd92 : y = 16'd24263;  // 92^0.7 ~= 23.694714
            8'd93 : y = 16'd24448;  // 93^0.7 ~= 23.874708
            8'd94 : y = 16'd24631;  // 94^0.7 ~= 24.054121
            8'd95 : y = 16'd24815;  // 95^0.7 ~= 24.232963
            8'd96 : y = 16'd24997;  // 96^0.7 ~= 24.411241
            8'd97 : y = 16'd25179;  // 97^0.7 ~= 24.588963
            8'd98 : y = 16'd25361;  // 98^0.7 ~= 24.766136
            8'd99 : y = 16'd25541;  // 99^0.7 ~= 24.942767
            8'd100: y = 16'd25722;  // 100^0.7 ~= 25.118864
            8'd101: y = 16'd25902;  // 101^0.7 ~= 25.294434
            8'd102: y = 16'd26081;  // 102^0.7 ~= 25.469482
            8'd103: y = 16'd26259;  // 103^0.7 ~= 25.644017
            8'd104: y = 16'd26438;  // 104^0.7 ~= 25.818044
            8'd105: y = 16'd26615;  // 105^0.7 ~= 25.991570
            8'd106: y = 16'd26793;  // 106^0.7 ~= 26.164600
            8'd107: y = 16'd26969;  // 107^0.7 ~= 26.337142
            8'd108: y = 16'd27145;  // 108^0.7 ~= 26.509200
            8'd109: y = 16'd27321;  // 109^0.7 ~= 26.680782
            8'd110: y = 16'd27496;  // 110^0.7 ~= 26.851891
            8'd111: y = 16'd27671;  // 111^0.7 ~= 27.022535
            8'd112: y = 16'd27845;  // 112^0.7 ~= 27.192718
            8'd113: y = 16'd28019;  // 113^0.7 ~= 27.362446
            8'd114: y = 16'd28192;  // 114^0.7 ~= 27.531723
            8'd115: y = 16'd28365;  // 115^0.7 ~= 27.700556
            8'd116: y = 16'd28538;  // 116^0.7 ~= 27.868949
            8'd117: y = 16'd28710;  // 117^0.7 ~= 28.036907
            8'd118: y = 16'd28881;  // 118^0.7 ~= 28.204435
            8'd119: y = 16'd29052;  // 119^0.7 ~= 28.371538
            8'd120: y = 16'd29223;  // 120^0.7 ~= 28.538219
            8'd121: y = 16'd29393;  // 121^0.7 ~= 28.704485
            8'd122: y = 16'd29563;  // 122^0.7 ~= 28.870339
            8'd123: y = 16'd29733;  // 123^0.7 ~= 29.035785
            8'd124: y = 16'd29902;  // 124^0.7 ~= 29.200829
            8'd125: y = 16'd30070;  // 125^0.7 ~= 29.365474
            8'd126: y = 16'd30238;  // 126^0.7 ~= 29.529724
            8'd127: y = 16'd30406;  // 127^0.7 ~= 29.693583
            8'd128: y = 16'd30574;  // 128^0.7 ~= 29.857056
            8'd129: y = 16'd30741;  // 129^0.7 ~= 30.020146
            8'd130: y = 16'd30907;  // 130^0.7 ~= 30.182857
            8'd131: y = 16'd31073;  // 131^0.7 ~= 30.345193
            8'd132: y = 16'd31239;  // 132^0.7 ~= 30.507158
            8'd133: y = 16'd31405;  // 133^0.7 ~= 30.668755
            8'd134: y = 16'd31570;  // 134^0.7 ~= 30.829988
            8'd135: y = 16'd31735;  // 135^0.7 ~= 30.990861
            8'd136: y = 16'd31899;  // 136^0.7 ~= 31.151376
            8'd137: y = 16'd32063;  // 137^0.7 ~= 31.311538
            8'd138: y = 16'd32227;  // 138^0.7 ~= 31.471349
            8'd139: y = 16'd32390;  // 139^0.7 ~= 31.630813
            8'd140: y = 16'd32553;  // 140^0.7 ~= 31.789934
            8'd141: y = 16'd32715;  // 141^0.7 ~= 31.948714
            8'd142: y = 16'd32878;  // 142^0.7 ~= 32.107156
            8'd143: y = 16'd33040;  // 143^0.7 ~= 32.265264
            8'd144: y = 16'd33201;  // 144^0.7 ~= 32.423041
            8'd145: y = 16'd33362;  // 145^0.7 ~= 32.580489
            8'd146: y = 16'd33523;  // 146^0.7 ~= 32.737612
            8'd147: y = 16'd33684;  // 147^0.7 ~= 32.894413
            8'd148: y = 16'd33844;  // 148^0.7 ~= 33.050893
            8'd149: y = 16'd34004;  // 149^0.7 ~= 33.207057
            8'd150: y = 16'd34164;  // 150^0.7 ~= 33.362907
            8'd151: y = 16'd34323;  // 151^0.7 ~= 33.518445
            8'd152: y = 16'd34482;  // 152^0.7 ~= 33.673675
            8'd153: y = 16'd34640;  // 153^0.7 ~= 33.828598
            8'd154: y = 16'd34799;  // 154^0.7 ~= 33.983218
            8'd155: y = 16'd34957;  // 155^0.7 ~= 34.137537
            8'd156: y = 16'd35115;  // 156^0.7 ~= 34.291558
            8'd157: y = 16'd35272;  // 157^0.7 ~= 34.445283
            8'd158: y = 16'd35429;  // 158^0.7 ~= 34.598714
            8'd159: y = 16'd35586;  // 159^0.7 ~= 34.751855
            8'd160: y = 16'd35742;  // 160^0.7 ~= 34.904706
            8'd161: y = 16'd35899;  // 161^0.7 ~= 35.057272
            8'd162: y = 16'd36055;  // 162^0.7 ~= 35.209553
            8'd163: y = 16'd36210;  // 163^0.7 ~= 35.361552
            8'd164: y = 16'd36366;  // 164^0.7 ~= 35.513272
            8'd165: y = 16'd36521;  // 165^0.7 ~= 35.664715
            8'd166: y = 16'd36675;  // 166^0.7 ~= 35.815883
            8'd167: y = 16'd36830;  // 167^0.7 ~= 35.966778
            8'd168: y = 16'd36984;  // 168^0.7 ~= 36.117402
            8'd169: y = 16'd37138;  // 169^0.7 ~= 36.267757
            8'd170: y = 16'd37292;  // 170^0.7 ~= 36.417845
            8'd171: y = 16'd37445;  // 171^0.7 ~= 36.567669
            8'd172: y = 16'd37598;  // 172^0.7 ~= 36.717230
            8'd173: y = 16'd37751;  // 173^0.7 ~= 36.866531
            8'd174: y = 16'd37904;  // 174^0.7 ~= 37.015573
            8'd175: y = 16'd38056;  // 175^0.7 ~= 37.164358
            8'd176: y = 16'd38208;  // 176^0.7 ~= 37.312888
            8'd177: y = 16'd38360;  // 177^0.7 ~= 37.461166
            8'd178: y = 16'd38512;  // 178^0.7 ~= 37.609192
            8'd179: y = 16'd38663;  // 179^0.7 ~= 37.756969
            8'd180: y = 16'd38814;  // 180^0.7 ~= 37.904498
            8'd181: y = 16'd38965;  // 181^0.7 ~= 38.051782
            8'd182: y = 16'd39116;  // 182^0.7 ~= 38.198822
            8'd183: y = 16'd39266;  // 183^0.7 ~= 38.345620
            8'd184: y = 16'd39416;  // 184^0.7 ~= 38.492177
            8'd185: y = 16'd39566;  // 185^0.7 ~= 38.638496
            8'd186: y = 16'd39715;  // 186^0.7 ~= 38.784577
            8'd187: y = 16'd39865;  // 187^0.7 ~= 38.930423
            8'd188: y = 16'd40014;  // 188^0.7 ~= 39.076035
            8'd189: y = 16'd40163;  // 189^0.7 ~= 39.221415
            8'd190: y = 16'd40311;  // 190^0.7 ~= 39.366565
            8'd191: y = 16'd40460;  // 191^0.7 ~= 39.511485
            8'd192: y = 16'd40608;  // 192^0.7 ~= 39.656178
            8'd193: y = 16'd40756;  // 193^0.7 ~= 39.800646
            8'd194: y = 16'd40904;  // 194^0.7 ~= 39.944888
            8'd195: y = 16'd41051;  // 195^0.7 ~= 40.088908
            8'd196: y = 16'd41198;  // 196^0.7 ~= 40.232707
            8'd197: y = 16'd41345;  // 197^0.7 ~= 40.376285
            8'd198: y = 16'd41492;  // 198^0.7 ~= 40.519645
            8'd199: y = 16'd41639;  // 199^0.7 ~= 40.662788
            8'd200: y = 16'd41785;  // 200^0.7 ~= 40.805715
            8'd201: y = 16'd41931;  // 201^0.7 ~= 40.948429
            8'd202: y = 16'd42077;  // 202^0.7 ~= 41.090929
            8'd203: y = 16'd42223;  // 203^0.7 ~= 41.233218
            8'd204: y = 16'd42368;  // 204^0.7 ~= 41.375296
            8'd205: y = 16'd42514;  // 205^0.7 ~= 41.517166
            8'd206: y = 16'd42659;  // 206^0.7 ~= 41.658829
            8'd207: y = 16'd42803;  // 207^0.7 ~= 41.800285
            8'd208: y = 16'd42948;  // 208^0.7 ~= 41.941536
            8'd209: y = 16'd43093;  // 209^0.7 ~= 42.082584
            8'd210: y = 16'd43237;  // 210^0.7 ~= 42.223430
            8'd211: y = 16'd43381;  // 211^0.7 ~= 42.364074
            8'd212: y = 16'd43525;  // 212^0.7 ~= 42.504519
            8'd213: y = 16'd43668;  // 213^0.7 ~= 42.644765
            8'd214: y = 16'd43812;  // 214^0.7 ~= 42.784813
            8'd215: y = 16'd43955;  // 215^0.7 ~= 42.924666
            8'd216: y = 16'd44098;  // 216^0.7 ~= 43.064323
            8'd217: y = 16'd44241;  // 217^0.7 ~= 43.203787
            8'd218: y = 16'd44383;  // 218^0.7 ~= 43.343058
            8'd219: y = 16'd44526;  // 219^0.7 ~= 43.482137
            8'd220: y = 16'd44668;  // 220^0.7 ~= 43.621026
            8'd221: y = 16'd44810;  // 221^0.7 ~= 43.759726
            8'd222: y = 16'd44952;  // 222^0.7 ~= 43.898237
            8'd223: y = 16'd45093;  // 223^0.7 ~= 44.036562
            8'd224: y = 16'd45235;  // 224^0.7 ~= 44.174700
            8'd225: y = 16'd45376;  // 225^0.7 ~= 44.312654
            8'd226: y = 16'd45517;  // 226^0.7 ~= 44.450424
            8'd227: y = 16'd45658;  // 227^0.7 ~= 44.588011
            8'd228: y = 16'd45799;  // 228^0.7 ~= 44.725416
            8'd229: y = 16'd45939;  // 229^0.7 ~= 44.862641
            8'd230: y = 16'd46080;  // 230^0.7 ~= 44.999686
            8'd231: y = 16'd46220;  // 231^0.7 ~= 45.136553
            8'd232: y = 16'd46360;  // 232^0.7 ~= 45.273241
            8'd233: y = 16'd46500;  // 233^0.7 ~= 45.409754
            8'd234: y = 16'd46639;  // 234^0.7 ~= 45.546090
            8'd235: y = 16'd46779;  // 235^0.7 ~= 45.682252
            8'd236: y = 16'd46918;  // 236^0.7 ~= 45.818240
            8'd237: y = 16'd47057;  // 237^0.7 ~= 45.954055
            8'd238: y = 16'd47196;  // 238^0.7 ~= 46.089699
            8'd239: y = 16'd47335;  // 239^0.7 ~= 46.225171
            8'd240: y = 16'd47473;  // 240^0.7 ~= 46.360474
            8'd241: y = 16'd47612;  // 241^0.7 ~= 46.495608
            8'd242: y = 16'd47750;  // 242^0.7 ~= 46.630573
            8'd243: y = 16'd47888;  // 243^0.7 ~= 46.765372
            8'd244: y = 16'd48026;  // 244^0.7 ~= 46.900004
            8'd245: y = 16'd48163;  // 245^0.7 ~= 47.034470
            8'd246: y = 16'd48301;  // 246^0.7 ~= 47.168773
            8'd247: y = 16'd48438;  // 247^0.7 ~= 47.302911
            8'd248: y = 16'd48575;  // 248^0.7 ~= 47.436887
            8'd249: y = 16'd48712;  // 249^0.7 ~= 47.570700
            8'd250: y = 16'd48849;  // 250^0.7 ~= 47.704353
            8'd251: y = 16'd48986;  // 251^0.7 ~= 47.837845
            8'd252: y = 16'd49122;  // 252^0.7 ~= 47.971177
            8'd253: y = 16'd49259;  // 253^0.7 ~= 48.104352
            8'd254: y = 16'd49395;  // 254^0.7 ~= 48.237368
            8'd255: y = 16'd49531;  // 255^0.7 ~= 48.370227
            default: y = 16'd0;
        endcase
    end
endmodule
