// Transmission Estimation, Scene Recovery and Saturation Correction Module
`define Image_Size (512 * 512)
module TE_and_SRSC (
    input        clk,
    input        rst,
    
    input        input_valid,                                 // Input data valid signal
    input [23:0] input_pixel_1, input_pixel_2, input_pixel_3,
                 input_pixel_4, input_pixel_5, input_pixel_6,
                 input_pixel_7, input_pixel_8, input_pixel_9, // 3x3 window input
    
    input  [7:0] A_R, A_G, A_B,                               // Atmospheric Light Values
    input [15:0] Inv_AR, Inv_AG, Inv_AB,                      // Inverse Atmospheric Light Values(Q0.16)

    output [7:0] J_R, J_G, J_B,                               // Output corrected pixels
    output       output_valid                                 // Output data valid signal
);

    // Pipeline the Center Pixel for SRSC
    reg [23:0] I_0_P, I_1_P, I_2_P;
    
    // Pipeline Atmospheric Light values for SRSC
    reg [7:0] A_R0_P, A_G0_P, A_B0_P;
    reg [7:0] A_R1_P, A_G1_P, A_B1_P;
    reg [7:0] A_R2_P, A_G2_P, A_B2_P;
    
    //==================================================================================
    // STAGE 4 LOGIC
    //==================================================================================
    
    // Detect the type of edge in the 3x3 window
    wire [1:0] ed1, ed2, ed3;
    
    // Pipeline Registers
    reg [1:0] window_edge_P;
    
    reg [15:0] Inv_AR_P, Inv_AG_P, Inv_AB_P;
    
    reg [23:0] I1_P, I2_P, I3_P,
               I4_P, I5_P, I6_P,
               I7_P, I8_P, I9_P;
               
    reg        stage_4_valid;
    
    //===========================================
    // Detect the type of edge in the 3x3 window
    ED_Top EdgeDetection (
        .input_pixel_1(input_pixel_1), .input_pixel_2(input_pixel_2), .input_pixel_3(input_pixel_3),
        .input_pixel_4(input_pixel_4),                                .input_pixel_6(input_pixel_6), 
        .input_pixel_7(input_pixel_7), .input_pixel_8(input_pixel_8), .input_pixel_9(input_pixel_9),
        
        .ED1_out(ed1), .ED2_out(ed2), .ED3_out(ed3)
    );
    //===========================================
    
    // Update Stage 4 Pipeline Registers
    always @(posedge clk) begin
        if (rst) begin
            window_edge_P <= 0;
        
            I1_P <= 0; I2_P <= 0; I3_P <= 0;
            I4_P <= 0; I5_P <= 0; I6_P <= 0;
            I7_P <= 0; I8_P <= 0; I9_P <= 0;
                
            Inv_AR_P <= 0; Inv_AG_P <= 0; Inv_AB_P <= 0;
                    
            I_0_P <= 0;
            A_R0_P <= 0; A_G0_P <= 0; A_B0_P <= 0;
                    
            stage_4_valid <= 0;
        end
        else begin
            window_edge_P <= (ed1 > ed2) ? ((ed1 > ed3) ? ed1 : ed3) : ((ed2 > ed3) ? ed2 : ed3);
        
            I1_P <= input_pixel_1; I2_P <= input_pixel_2; I3_P <= input_pixel_3;
            I4_P <= input_pixel_4; I5_P <= input_pixel_5; I6_P <= input_pixel_6;
            I7_P <= input_pixel_7; I8_P <= input_pixel_8; I9_P <= input_pixel_9;
                    
            Inv_AR_P <= Inv_AR; Inv_AG_P <= Inv_AG; Inv_AB_P <= Inv_AB;

            I_0_P <= input_pixel_5;
            A_R0_P <= A_R; A_G0_P <= A_G; A_B0_P <= A_B;
                    
            stage_4_valid <= input_valid;
        end
    end
    
    //==================================================================================
    // STAGE 5 LOGIC
    //==================================================================================
    
    // ? = 63/64
    parameter OMEGA_D = 4;
    
    wire [7:0] filtered_pixel_red, filtered_pixel_green, filtered_pixel_blue;
    
    // Pipeline Registers
    reg [15:0] Inv_AR_P1, Inv_AG_P1, Inv_AB_P1;
    
    reg [7:0] filtered_pixel_red_P, filtered_pixel_green_P, filtered_pixel_blue_P;
    
    reg stage_5_valid;
    
    //===========================================
    // Filter blocks to apply Gaussian Filter or Mean Filter based on the edge detected
    WindowFilter Red_WindowFilter (
        .window_edge(window_edge_P),
    
        .input_pixel_1(I1_P[23:16]), .input_pixel_2(I2_P[23:16]), .input_pixel_3(I3_P[23:16]),
        .input_pixel_4(I4_P[23:16]), .input_pixel_5(I5_P[23:16]), .input_pixel_6(I6_P[23:16]),
        .input_pixel_7(I7_P[23:16]), .input_pixel_8(I8_P[23:16]), .input_pixel_9(I9_P[23:16]),
        
        .filtered_pixel(filtered_pixel_red)
    );
                   
    WindowFilter Green_WindowFilter (
        .window_edge(window_edge_P),

        .input_pixel_1(I1_P[15:8]), .input_pixel_2(I2_P[15:8]), .input_pixel_3(I3_P[15:8]),
        .input_pixel_4(I4_P[15:8]), .input_pixel_5(I5_P[15:8]), .input_pixel_6(I6_P[15:8]),
        .input_pixel_7(I7_P[15:8]), .input_pixel_8(I8_P[15:8]), .input_pixel_9(I9_P[15:8]),
        
        .filtered_pixel(filtered_pixel_green)
    );
                   
    WindowFilter Blue_WindowFilter (
        .window_edge(window_edge_P),

        .input_pixel_1(I1_P[7:0]), .input_pixel_2(I2_P[7:0]), .input_pixel_3(I3_P[7:0]),
        .input_pixel_4(I4_P[7:0]), .input_pixel_5(I5_P[7:0]), .input_pixel_6(I6_P[7:0]),
        .input_pixel_7(I7_P[7:0]), .input_pixel_8(I8_P[7:0]), .input_pixel_9(I9_P[7:0]),
                       
        .filtered_pixel(filtered_pixel_blue)
    );
    //===========================================
    
    // Update Stage 5 Pipeline Registers 
    always @(posedge clk) begin
        if (rst) begin
            
            Inv_AR_P1 <= 0; Inv_AG_P1 <= 0; Inv_AB_P1 <= 0;
            
            filtered_pixel_red_P <= 0; filtered_pixel_green_P <= 0; filtered_pixel_blue_P <= 0;
            
            I_1_P <= 0;
            A_R1_P <= 0; A_G1_P <= 0; A_B1_P <= 0;
            
            stage_5_valid <= 0;
        end
        else begin
            // Apply the scaling factor ? = 63/64 to the Inverse Atmospheric Light values
            Inv_AR_P1 <= Inv_AR_P - (Inv_AR_P >> OMEGA_D);
            Inv_AG_P1 <= Inv_AG_P - (Inv_AG_P >> OMEGA_D);
            Inv_AB_P1 <= Inv_AB_P - (Inv_AB_P >> OMEGA_D);
            
            filtered_pixel_red_P <= filtered_pixel_red;
            filtered_pixel_green_P <= filtered_pixel_green;
            filtered_pixel_blue_P <= filtered_pixel_blue;
                                
            I_1_P <= I_0_P;
                                
            A_R1_P <= A_R0_P; A_G1_P <= A_G0_P; A_B1_P <= A_B0_P;
                                
            stage_5_valid <= stage_4_valid;
        end
    end
    
    //==========================================================================
    // STAGE 6 LOGIC
    //==========================================================================
    
    // Select signal for minimum filter result
    wire  [1:0] min_val_sel;
    
    wire [7:0] min_Fc;
    
    wire [15:0] min_Ac;
        
    wire [13:0] product;
    
    reg         stage_6_valid;
    
    //===========================================
    // Comparator to determine the minimum value of the filter results
    Comparator_Minimum Minimum_Filter_Select (
        .red(filtered_pixel_red_P), .green(filtered_pixel_green_P), .blue(filtered_pixel_blue_P),
        
        .min_val_sel(min_val_sel)
    );
    
    // Multiplexer to choose minimum of the filter results
    Filter_Result_Multiplexer Minimum_Filtered_Pixel_Result (
        .F_R(filtered_pixel_red_P), .F_G(filtered_pixel_green_P), .F_B(filtered_pixel_blue_P),
        
        .sel(min_val_sel),
        
        .Fc(min_Fc)
    );
    
    // Multiplexer to choose minimum of Atmospheric Light values
    Inv_Ac_Multiplexer Minimum_Inv_ALE_Value (
        .Inv_AR(Inv_AR_P1), .Inv_AG(Inv_AG_P1), .Inv_AB(Inv_AB_P1),
        
        .sel(min_val_sel),
        
        .Inv_Ac(min_Ac)
    );
    
    // Multiplier modules to compute Fc * ?/Ac
    Multiplier_TE Fc_InvAc_Multiplier (
        .clk(clk), .rst(rst),
        
        .Fc(min_Fc),
        .Inv_Ac(min_Ac),
        
        .product(product)
    );
    //===========================================
    
    // Update Stage 6 Pipeline Registers
    always @(posedge clk) begin
        if (rst) begin
            I_2_P <= 0;
            A_R2_P <= 0; A_G2_P <= 0; A_B2_P <= 0;
            
            stage_6_valid <= 0;
        end
        else begin
            I_2_P <= I_1_P;
            A_R2_P <= A_R1_P; A_G2_P <= A_G1_P; A_B2_P <= A_B1_P;
            
            stage_6_valid <= stage_5_valid;
        end
    end
    
    //==========================================================================
    // STAGE 7 LOGIC
    //==========================================================================
    // Transmission value in Q0.14
    wire [13:0] transmission;
    
    // Compute (|Ic - Ac|)
    wire [7:0]  IR_minus_AR, IG_minus_AG, IB_minus_AB;
    wire        add_or_sub_R, add_or_sub_G, add_or_sub_B;
    wire [7:0] I_R = I_2_P[23:16], I_G = I_2_P[15:8], I_B = I_2_P[7:0];
    
    // Pipeline Registers for stage 7
    reg [13:0]  transmission_P;
    
    reg [7:0]   A_R_P, A_G_P, A_B_P;
    reg [7:0]   I_R_P, I_G_P, I_B_P;
    
    reg [7:0]   IR_minus_AR_P, IG_minus_AG_P, IB_minus_AB_P;
    reg         add_or_sub_R_P, add_or_sub_G_P, add_or_sub_B_P;
    
    reg         stage_7_valid;
    
    //===========================================
            
    // Subtractor to compute final transmission value
    Subtractor_TE Subtractor_TE (
        .in(product),
        .out(transmission)
    );
    
    // SUBTRACTOR MODULES TO COMPUTE (|Ic - Ac|)
    Subtractor_SRSC Sub_Red (
        .Ic(I_R),
        .Ac(A_R2_P),
        
        .diff(IR_minus_AR),
        
        .add_or_sub(add_or_sub_R)
    );
                
    Subtractor_SRSC Sub_Green (
        .Ic(I_G),
        .Ac(A_G2_P),
        
        .diff(IG_minus_AG),
        
        .add_or_sub(add_or_sub_G)
    );
            
    Subtractor_SRSC Sub_Blue (
        .Ic(I_B),
        .Ac(A_B2_P),
        
        .diff(IB_minus_AB),
        
        .add_or_sub(add_or_sub_B)
    );
    //===========================================
    
    // Update Stage 7 Pipeline Registers
    always @(posedge clk) begin
        if (rst) begin
            transmission_P <= 0;
            
            A_R_P <= 0;
            A_G_P <= 0;
            A_B_P <= 0;
            
            I_R_P <= 0;
            I_G_P <= 0;
            I_B_P <= 0;
            
            IR_minus_AR_P <= 0;
            IG_minus_AG_P <= 0;
            IB_minus_AB_P <= 0;
            
            add_or_sub_R_P <= 0;
            add_or_sub_G_P <= 0;
            add_or_sub_B_P <= 0;
            
            stage_7_valid <= 0;
        end
        else begin
            transmission_P <= transmission;
            
            A_R_P <= A_R2_P;
            A_G_P <= A_G2_P;
            A_B_P <= A_B2_P;
            
            I_R_P <= I_R;
            I_G_P <= I_G;
            I_B_P <= I_B;
            
            IR_minus_AR_P <= IR_minus_AR;
            IG_minus_AG_P <= IG_minus_AG;
            IB_minus_AB_P <= IB_minus_AB;
            
            add_or_sub_R_P <= add_or_sub_R;
            add_or_sub_G_P <= add_or_sub_G;
            add_or_sub_B_P <= add_or_sub_B;
            
            stage_7_valid <= stage_6_valid;
        end
    end
                
    //==========================================================================
    // STAGE 8 LOGIC
    //==========================================================================
                
    wire [13:0] inverse_transmission;

    // Compute (|Ic-Ac|)*(1/T)
    wire [7:0]  IR_minus_AR_x_T, IG_minus_AG_x_T, IB_minus_AB_x_T;

    // Pipeline Registers for stage 8
    reg [7:0]   A_R_P1, A_G_P1, A_B_P1;
    reg [7:0]   I_R_P1, I_G_P1, I_B_P1;
    
    reg         add_or_sub_R_P1, add_or_sub_G_P1, add_or_sub_B_P1;
    
    reg         stage_8_valid;
    
    //===========================================
    // TRANSMISSION RECIPROCAL LOOKUP TABLE
    Transmission_Reciprocal_LUT Transmission_Reciprocal_LUT (
        .in(transmission_P),
                        
        .out(inverse_transmission)
    );
                
    // MULTIPLIER MODULES TO COMPUTE (|Ic-Ac|)*(1/T)
    Multiplier_SRSC Mult_Red (
        .clk(clk), .rst(rst),
        
        .Inv_Trans(inverse_transmission),
        .Ic_minus_Ac(IR_minus_AR_P),
        
        .result(IR_minus_AR_x_T)
    );
                        
    Multiplier_SRSC Mult_Green (
        .clk(clk), .rst(rst),
        
        .Inv_Trans(inverse_transmission),
        .Ic_minus_Ac(IG_minus_AG_P),
        
        .result(IG_minus_AG_x_T)
    );
                    
    Multiplier_SRSC Mult_Blue (
        .clk(clk), .rst(rst),
        
        .Inv_Trans(inverse_transmission),
        .Ic_minus_Ac(IB_minus_AB_P),
        
        .result(IB_minus_AB_x_T)
    );
    //===========================================
    
    // Update stage 8 pipeline registers
    always @(posedge clk) begin
        if (rst) begin        
            A_R_P1 <= 0;
            A_G_P1 <= 0;
            A_B_P1 <= 0;
            
            I_R_P1 <= 0;
            I_G_P1 <= 0;
            I_B_P1 <= 0;
            
            add_or_sub_R_P1 <= 0;
            add_or_sub_G_P1 <= 0;
            add_or_sub_B_P1 <= 0;
            
            stage_8_valid <= 0;
        end
        else begin       
            A_R_P1 <= A_R_P;
            A_G_P1 <= A_G_P;
            A_B_P1 <= A_B_P;
            
            I_R_P1 <= I_R_P;
            I_G_P1 <= I_G_P;
            I_B_P1 <= I_B_P;
            
            add_or_sub_R_P1 <= add_or_sub_R_P;
            add_or_sub_G_P1 <= add_or_sub_G_P;
            add_or_sub_B_P1 <= add_or_sub_B_P;
            
            stage_8_valid <= stage_7_valid;
        end
    end
    
    //==========================================================================
    // STAGE 9 LOGIC
    //==========================================================================
    
    // Pipeline Registers for stage 9
    reg [7:0]  A_R_P2, A_G_P2, A_B_P2;
    reg [7:0]  I_R_P2, I_G_P2, I_B_P2;
    reg [7:0]  Mult_Red_P, Mult_Green_P, Mult_Blue_P;
    
    reg        add_or_sub_R_P2, add_or_sub_G_P2, add_or_sub_B_P2;
    
    reg        stage_9_valid;
    
    // Update stage 9 pipeline registers
    always @(posedge clk) begin
        if (rst) begin
            A_R_P2 <= 0;
            A_G_P2 <= 0;
            A_B_P2 <= 0;
            
            I_R_P2 <= 0;
            I_G_P2 <= 0;
            I_B_P2 <= 0;
            
            add_or_sub_R_P2 <= 0;
            add_or_sub_G_P2 <= 0;
            add_or_sub_B_P2 <= 0;
            
            Mult_Red_P <= 0;
            Mult_Green_P <= 0;
            Mult_Blue_P <= 0;
            
            stage_9_valid <= 0;
        end
        else begin
            A_R_P2 <= A_R_P1;
            A_G_P2 <= A_G_P1;
            A_B_P2 <= A_B_P1;
            
            I_R_P2 <= I_R_P1;
            I_G_P2 <= I_G_P1;
            I_B_P2 <= I_B_P1;
            
            add_or_sub_R_P2 <= add_or_sub_R_P1;
            add_or_sub_G_P2 <= add_or_sub_G_P1;
            add_or_sub_B_P2 <= add_or_sub_B_P1;
            
            Mult_Red_P <= IR_minus_AR_x_T;
            Mult_Green_P <= IG_minus_AG_x_T;
            Mult_Blue_P <= IB_minus_AB_x_T;
            
            stage_9_valid <= stage_8_valid;
        end
    end
    
    //==========================================================================
    // STAGE 10 LOGIC
    //==========================================================================
    
    // Compute Ac +/- (|Ic-Ac|/T)
    wire [7:0] Sum_Red, Sum_Green, Sum_Blue;
    
    // Outputs of Look-Up Tables for Saturation Corection
    wire [11:0] J_R_Corrected, J_G_Corrected, J_B_Corrected;
    wire [11:0] A_R_Corrected, A_G_Corrected, A_B_Corrected;

    // Pipeline Registers for stage 10
    reg       stage_10_valid;
    
    //===========================================
    // ADDER BLOCKS TO COMPUTE Ac +/- (|Ic-Ac|/T)
    Adder_SRSC Add_Red (
        .Ac(A_R_P2),
        .Ic(I_R_P2),
        .Multiplier_out(Mult_Red_P),
         
        .add_or_sub(add_or_sub_R_P2),
         
        .out(Sum_Red)
    );
                         
    Adder_SRSC Add_Green (
        .Ac(A_G_P2),
        .Ic(I_G_P2),
        .Multiplier_out(Mult_Green_P),
         
        .add_or_sub(add_or_sub_G_P2),
         
        .out(Sum_Green)
    );
                         
    Adder_SRSC Add_Blue (
        .Ac(A_B_P2),
        .Ic(I_B_P2),
        .Multiplier_out(Mult_Blue_P),
         
        .add_or_sub(add_or_sub_B_P2),
         
        .out(Sum_Blue)
    );
    
    // LOOK-UP TABLES TO COMPUTE Ac ^ ? AND Jc ^ (1 - ?) (? = 0.3)
    LUT_03 A_R_Correction (
        .in(A_R_P2),
        .out(A_R_Corrected)
    );
    
    LUT_03 A_G_Correction (
        .in(A_G_P2),
        .out(A_G_Corrected)
    );
    
    LUT_03 A_B_Correction (
        .in(A_B_P2),
        .out(A_B_Corrected)
    );
    
    LUT_07 J_R_Correction (
        .in(Sum_Red),
        .out(J_R_Corrected)
    );
    
    LUT_07 J_G_Correction (
        .in(Sum_Green),
        .out(J_G_Corrected)
    );
    
    LUT_07 J_B_Correction (
        .in(Sum_Blue),
        .out(J_B_Corrected)
    );
                    
    // MULTIPLIER MODULES TO COMPUTE Ac^? * Jc^(1-?)
    Saturation_Correction_Multiplier Saturation_Correction_Red (
        .clk(clk), .rst(rst),
        
        .x1(A_R_Corrected), .x2(J_R_Corrected),
        
        .result(J_R)
    );
    
    Saturation_Correction_Multiplier Saturation_Correction_Green (
        .clk(clk), .rst(rst),
        
        .x1(A_G_Corrected), .x2(J_G_Corrected),
        
        .result(J_G)
    );
    
    Saturation_Correction_Multiplier Saturation_Correction_Blue (
        .clk(clk), .rst(rst),
        
        .x1(A_B_Corrected), .x2(J_B_Corrected),
        
        .result(J_B)
    );
    //===========================================
    
    // Update stage 10 pipeline registers
    always @(posedge clk) begin
        if (rst) begin
            stage_10_valid <= 0;
        end
        else begin
            stage_10_valid <= stage_9_valid;
        end
    end

    // Stage 11 assignments
    assign output_valid = stage_10_valid;

endmodule
