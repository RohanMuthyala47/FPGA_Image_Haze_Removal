//module test(
//    input clk,
//    input rst,
//    input input_is_valid,

//    input wire [23:0] output_pixel_1,
//    input wire [23:0] output_pixel_2,
//    input wire [23:0] output_pixel_3,
//    input wire [23:0] output_pixel_4,
//    input wire [23:0] output_pixel_5,
//    input wire [23:0] output_pixel_6,
//    input wire [23:0] output_pixel_7,
//    input wire [23:0] output_pixel_8,
//    input wire [23:0] output_pixel_9,
    
//    output wire [23:0] out_pixel,
//    output wire output_is_valid
//);
//    assign out_pixel = output_pixel_5;
//    assign output_is_valid = input_is_valid;
//endmodule