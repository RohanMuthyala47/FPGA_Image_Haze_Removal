module Transmission_Reciprocal_LUT (
    input      [13:0] in,  // Q0.14 input (unsigned)
    output reg [13:0] out  // Q2.12 reciprocal output (unsigned)
);

    always @(*) begin
        if(in < 'd4096)
             out <= 14'h3FFF;
        else begin
        casez(in)
            14'd 4097: out = 14'h3FFC;
            14'd 4098: out = 14'h3FF8;
            14'd 4099: out = 14'h3FF4;
            14'd 4100: out = 14'h3FF0;
            14'd 4101: out = 14'h3FEC;
            14'd 4102: out = 14'h3FE8;
            14'd 4103: out = 14'h3FE4;
            14'd 4104: out = 14'h3FE0;
            14'd 4105: out = 14'h3FDC;
            14'd 4106: out = 14'h3FD8;
            14'd 4107: out = 14'h3FD4;
            14'd 4108: out = 14'h3FD0;
            14'd 4109: out = 14'h3FCC;
            14'd 4110: out = 14'h3FC8;
            14'd 4111: out = 14'h3FC4;
            14'd 4112: out = 14'h3FC0;
            14'd 4113: out = 14'h3FBC;
            14'd 4114: out = 14'h3FB8;
            14'd 4115: out = 14'h3FB4;
            14'd 4116: out = 14'h3FB0;
            14'd 4117: out = 14'h3FAC;
            14'd 4118: out = 14'h3FA8;
            14'd 4119: out = 14'h3FA5;
            14'd 4120: out = 14'h3FA1;
            14'd 4121: out = 14'h3F9D;
            14'd 4122: out = 14'h3F99;
            14'd 4123: out = 14'h3F95;
            14'd 4124: out = 14'h3F91;
            14'd 4125: out = 14'h3F8D;
            14'd 4126: out = 14'h3F89;
            14'd 4127: out = 14'h3F85;
            14'd 4128: out = 14'h3F81;
            14'd 4129: out = 14'h3F7D;
            14'd 4130: out = 14'h3F79;
            14'd 4131: out = 14'h3F75;
            14'd 4132: out = 14'h3F71;
            14'd 4133: out = 14'h3F6D;
            14'd 4134: out = 14'h3F69;
            14'd 4135: out = 14'h3F65;
            14'd 4136: out = 14'h3F62;
            14'd 4137: out = 14'h3F5E;
            14'd 4138: out = 14'h3F5A;
            14'd 4139: out = 14'h3F56;
            14'd 4140: out = 14'h3F52;
            14'd 4141: out = 14'h3F4E;
            14'd 4142: out = 14'h3F4A;
            14'd 4143: out = 14'h3F46;
            14'd 4144: out = 14'h3F42;
            14'd 4145: out = 14'h3F3E;
            14'd 4146: out = 14'h3F3A;
            14'd 4147: out = 14'h3F37;
            14'd 4148: out = 14'h3F33;
            14'd 4149: out = 14'h3F2F;
            14'd 4150: out = 14'h3F2B;
            14'd 4151: out = 14'h3F27;
            14'd 4152: out = 14'h3F23;
            14'd 4153: out = 14'h3F1F;
            14'd 4154: out = 14'h3F1B;
            14'd 4155: out = 14'h3F17;
            14'd 4156: out = 14'h3F13;
            14'd 4157: out = 14'h3F10;
            14'd 4158: out = 14'h3F0C;
            14'd 4159: out = 14'h3F08;
            14'd 4160: out = 14'h3F04;
            14'd 4161: out = 14'h3F00;
            14'd 4162: out = 14'h3EFC;
            14'd 4163: out = 14'h3EF8;
            14'd 4164: out = 14'h3EF4;
            14'd 4165: out = 14'h3EF1;
            14'd 4166: out = 14'h3EED;
            14'd 4167: out = 14'h3EE9;
            14'd 4168: out = 14'h3EE5;
            14'd 4169: out = 14'h3EE1;
            14'd 4170: out = 14'h3EDD;
            14'd 4171: out = 14'h3ED9;
            14'd 4172: out = 14'h3ED6;
            14'd 4173: out = 14'h3ED2;
            14'd 4174: out = 14'h3ECE;
            14'd 4175: out = 14'h3ECA;
            14'd 4176: out = 14'h3EC6;
            14'd 4177: out = 14'h3EC2;
            14'd 4178: out = 14'h3EBE;
            14'd 4179: out = 14'h3EBB;
            14'd 4180: out = 14'h3EB7;
            14'd 4181: out = 14'h3EB3;
            14'd 4182: out = 14'h3EAF;
            14'd 4183: out = 14'h3EAB;
            14'd 4184: out = 14'h3EA7;
            14'd 4185: out = 14'h3EA4;
            14'd 4186: out = 14'h3EA0;
            14'd 4187: out = 14'h3E9C;
            14'd 4188: out = 14'h3E98;
            14'd 4189: out = 14'h3E94;
            14'd 4190: out = 14'h3E90;
            14'd 4191: out = 14'h3E8D;
            14'd 4192: out = 14'h3E89;
            14'd 4193: out = 14'h3E85;
            14'd 4194: out = 14'h3E81;
            14'd 4195: out = 14'h3E7D;
            14'd 4196: out = 14'h3E7A;
            14'd 4197: out = 14'h3E76;
            14'd 4198: out = 14'h3E72;
            14'd 4199: out = 14'h3E6E;
            14'd 4200: out = 14'h3E6A;
            14'd 4201: out = 14'h3E66;
            14'd 4202: out = 14'h3E63;
            14'd 4203: out = 14'h3E5F;
            14'd 4204: out = 14'h3E5B;
            14'd 4205: out = 14'h3E57;
            14'd 4206: out = 14'h3E54;
            14'd 4207: out = 14'h3E50;
            14'd 4208: out = 14'h3E4C;
            14'd 4209: out = 14'h3E48;
            14'd 4210: out = 14'h3E44;
            14'd 4211: out = 14'h3E41;
            14'd 4212: out = 14'h3E3D;
            14'd 4213: out = 14'h3E39;
            14'd 4214: out = 14'h3E35;
            14'd 4215: out = 14'h3E31;
            14'd 4216: out = 14'h3E2E;
            14'd 4217: out = 14'h3E2A;
            14'd 4218: out = 14'h3E26;
            14'd 4219: out = 14'h3E22;
            14'd 4220: out = 14'h3E1F;
            14'd 4221: out = 14'h3E1B;
            14'd 4222: out = 14'h3E17;
            14'd 4223: out = 14'h3E13;
            14'd 4224: out = 14'h3E10;
            14'd 4225: out = 14'h3E0C;
            14'd 4226: out = 14'h3E08;
            14'd 4227: out = 14'h3E04;
            14'd 4228: out = 14'h3E00;
            14'd 4229: out = 14'h3DFD;
            14'd 4230: out = 14'h3DF9;
            14'd 4231: out = 14'h3DF5;
            14'd 4232: out = 14'h3DF1;
            14'd 4233: out = 14'h3DEE;
            14'd 4234: out = 14'h3DEA;
            14'd 4235: out = 14'h3DE6;
            14'd 4236: out = 14'h3DE3;
            14'd 4237: out = 14'h3DDF;
            14'd 4238: out = 14'h3DDB;
            14'd 4239: out = 14'h3DD7;
            14'd 4240: out = 14'h3DD4;
            14'd 4241: out = 14'h3DD0;
            14'd 4242: out = 14'h3DCC;
            14'd 4243: out = 14'h3DC8;
            14'd 4244: out = 14'h3DC5;
            14'd 4245: out = 14'h3DC1;
            14'd 4246: out = 14'h3DBD;
            14'd 4247: out = 14'h3DB9;
            14'd 4248: out = 14'h3DB6;
            14'd 4249: out = 14'h3DB2;
            14'd 4250: out = 14'h3DAE;
            14'd 4251: out = 14'h3DAB;
            14'd 4252: out = 14'h3DA7;
            14'd 4253: out = 14'h3DA3;
            14'd 4254: out = 14'h3D9F;
            14'd 4255: out = 14'h3D9C;
            14'd 4256: out = 14'h3D98;
            14'd 4257: out = 14'h3D94;
            14'd 4258: out = 14'h3D91;
            14'd 4259: out = 14'h3D8D;
            14'd 4260: out = 14'h3D89;
            14'd 4261: out = 14'h3D86;
            14'd 4262: out = 14'h3D82;
            14'd 4263: out = 14'h3D7E;
            14'd 4264: out = 14'h3D7A;
            14'd 4265: out = 14'h3D77;
            14'd 4266: out = 14'h3D73;
            14'd 4267: out = 14'h3D6F;
            14'd 4268: out = 14'h3D6C;
            14'd 4269: out = 14'h3D68;
            14'd 4270: out = 14'h3D64;
            14'd 4271: out = 14'h3D61;
            14'd 4272: out = 14'h3D5D;
            14'd 4273: out = 14'h3D59;
            14'd 4274: out = 14'h3D56;
            14'd 4275: out = 14'h3D52;
            14'd 4276: out = 14'h3D4E;
            14'd 4277: out = 14'h3D4B;
            14'd 4278: out = 14'h3D47;
            14'd 4279: out = 14'h3D43;
            14'd 4280: out = 14'h3D40;
            14'd 4281: out = 14'h3D3C;
            14'd 4282: out = 14'h3D38;
            14'd 4283: out = 14'h3D35;
            14'd 4284: out = 14'h3D31;
            14'd 4285: out = 14'h3D2D;
            14'd 4286: out = 14'h3D2A;
            14'd 4287: out = 14'h3D26;
            14'd 4288: out = 14'h3D22;
            14'd 4289: out = 14'h3D1F;
            14'd 4290: out = 14'h3D1B;
            14'd 4291: out = 14'h3D17;
            14'd 4292: out = 14'h3D14;
            14'd 4293: out = 14'h3D10;
            14'd 4294: out = 14'h3D0D;
            14'd 4295: out = 14'h3D09;
            14'd 4296: out = 14'h3D05;
            14'd 4297: out = 14'h3D02;
            14'd 4298: out = 14'h3CFE;
            14'd 4299: out = 14'h3CFA;
            14'd 4300: out = 14'h3CF7;
            14'd 4301: out = 14'h3CF3;
            14'd 4302: out = 14'h3CEF;
            14'd 4303: out = 14'h3CEC;
            14'd 4304: out = 14'h3CE8;
            14'd 4305: out = 14'h3CE5;
            14'd 4306: out = 14'h3CE1;
            14'd 4307: out = 14'h3CDD;
            14'd 4308: out = 14'h3CDA;
            14'd 4309: out = 14'h3CD6;
            14'd 4310: out = 14'h3CD3;
            14'd 4311: out = 14'h3CCF;
            14'd 4312: out = 14'h3CCB;
            14'd 4313: out = 14'h3CC8;
            14'd 4314: out = 14'h3CC4;
            14'd 4315: out = 14'h3CC0;
            14'd 4316: out = 14'h3CBD;
            14'd 4317: out = 14'h3CB9;
            14'd 4318: out = 14'h3CB6;
            14'd 4319: out = 14'h3CB2;
            14'd 4320: out = 14'h3CAE;
            14'd 4321: out = 14'h3CAB;
            14'd 4322: out = 14'h3CA7;
            14'd 4323: out = 14'h3CA4;
            14'd 4324: out = 14'h3CA0;
            14'd 4325: out = 14'h3C9D;
            14'd 4326: out = 14'h3C99;
            14'd 4327: out = 14'h3C95;
            14'd 4328: out = 14'h3C92;
            14'd 4329: out = 14'h3C8E;
            14'd 4330: out = 14'h3C8B;
            14'd 4331: out = 14'h3C87;
            14'd 4332: out = 14'h3C83;
            14'd 4333: out = 14'h3C80;
            14'd 4334: out = 14'h3C7C;
            14'd 4335: out = 14'h3C79;
            14'd 4336: out = 14'h3C75;
            14'd 4337: out = 14'h3C72;
            14'd 4338: out = 14'h3C6E;
            14'd 4339: out = 14'h3C6A;
            14'd 4340: out = 14'h3C67;
            14'd 4341: out = 14'h3C63;
            14'd 4342: out = 14'h3C60;
            14'd 4343: out = 14'h3C5C;
            14'd 4344: out = 14'h3C59;
            14'd 4345: out = 14'h3C55;
            14'd 4346: out = 14'h3C52;
            14'd 4347: out = 14'h3C4E;
            14'd 4348: out = 14'h3C4A;
            14'd 4349: out = 14'h3C47;
            14'd 4350: out = 14'h3C43;
            14'd 4351: out = 14'h3C40;
            14'd 4352: out = 14'h3C3C;
            14'd 4353: out = 14'h3C39;
            14'd 4354: out = 14'h3C35;
            14'd 4355: out = 14'h3C32;
            14'd 4356: out = 14'h3C2E;
            14'd 4357: out = 14'h3C2B;
            14'd 4358: out = 14'h3C27;
            14'd 4359: out = 14'h3C23;
            14'd 4360: out = 14'h3C20;
            14'd 4361: out = 14'h3C1C;
            14'd 4362: out = 14'h3C19;
            14'd 4363: out = 14'h3C15;
            14'd 4364: out = 14'h3C12;
            14'd 4365: out = 14'h3C0E;
            14'd 4366: out = 14'h3C0B;
            14'd 4367: out = 14'h3C07;
            14'd 4368: out = 14'h3C04;
            14'd 4369: out = 14'h3C00;
            14'd 4370: out = 14'h3BFD;
            14'd 4371: out = 14'h3BF9;
            14'd 4372: out = 14'h3BF6;
            14'd 4373: out = 14'h3BF2;
            14'd 4374: out = 14'h3BEF;
            14'd 4375: out = 14'h3BEB;
            14'd 4376: out = 14'h3BE8;
            14'd 4377: out = 14'h3BE4;
            14'd 4378: out = 14'h3BE1;
            14'd 4379: out = 14'h3BDD;
            14'd 4380: out = 14'h3BDA;
            14'd 4381: out = 14'h3BD6;
            14'd 4382: out = 14'h3BD3;
            14'd 4383: out = 14'h3BCF;
            14'd 4384: out = 14'h3BCC;
            14'd 4385: out = 14'h3BC8;
            14'd 4386: out = 14'h3BC5;
            14'd 4387: out = 14'h3BC1;
            14'd 4388: out = 14'h3BBE;
            14'd 4389: out = 14'h3BBA;
            14'd 4390: out = 14'h3BB7;
            14'd 4391: out = 14'h3BB3;
            14'd 4392: out = 14'h3BB0;
            14'd 4393: out = 14'h3BAC;
            14'd 4394: out = 14'h3BA9;
            14'd 4395: out = 14'h3BA5;
            14'd 4396: out = 14'h3BA2;
            14'd 4397: out = 14'h3B9E;
            14'd 4398: out = 14'h3B9B;
            14'd 4399: out = 14'h3B97;
            14'd 4400: out = 14'h3B94;
            14'd 4401: out = 14'h3B91;
            14'd 4402: out = 14'h3B8D;
            14'd 4403: out = 14'h3B8A;
            14'd 4404: out = 14'h3B86;
            14'd 4405: out = 14'h3B83;
            14'd 4406: out = 14'h3B7F;
            14'd 4407: out = 14'h3B7C;
            14'd 4408: out = 14'h3B78;
            14'd 4409: out = 14'h3B75;
            14'd 4410: out = 14'h3B71;
            14'd 4411: out = 14'h3B6E;
            14'd 4412: out = 14'h3B6B;
            14'd 4413: out = 14'h3B67;
            14'd 4414: out = 14'h3B64;
            14'd 4415: out = 14'h3B60;
            14'd 4416: out = 14'h3B5D;
            14'd 4417: out = 14'h3B59;
            14'd 4418: out = 14'h3B56;
            14'd 4419: out = 14'h3B52;
            14'd 4420: out = 14'h3B4F;
            14'd 4421: out = 14'h3B4C;
            14'd 4422: out = 14'h3B48;
            14'd 4423: out = 14'h3B45;
            14'd 4424: out = 14'h3B41;
            14'd 4425: out = 14'h3B3E;
            14'd 4426: out = 14'h3B3A;
            14'd 4427: out = 14'h3B37;
            14'd 4428: out = 14'h3B34;
            14'd 4429: out = 14'h3B30;
            14'd 4430: out = 14'h3B2D;
            14'd 4431: out = 14'h3B29;
            14'd 4432: out = 14'h3B26;
            14'd 4433: out = 14'h3B22;
            14'd 4434: out = 14'h3B1F;
            14'd 4435: out = 14'h3B1C;
            14'd 4436: out = 14'h3B18;
            14'd 4437: out = 14'h3B15;
            14'd 4438: out = 14'h3B11;
            14'd 4439: out = 14'h3B0E;
            14'd 4440: out = 14'h3B0B;
            14'd 4441: out = 14'h3B07;
            14'd 4442: out = 14'h3B04;
            14'd 4443: out = 14'h3B00;
            14'd 4444: out = 14'h3AFD;
            14'd 4445: out = 14'h3AFA;
            14'd 4446: out = 14'h3AF6;
            14'd 4447: out = 14'h3AF3;
            14'd 4448: out = 14'h3AEF;
            14'd 4449: out = 14'h3AEC;
            14'd 4450: out = 14'h3AE9;
            14'd 4451: out = 14'h3AE5;
            14'd 4452: out = 14'h3AE2;
            14'd 4453: out = 14'h3ADE;
            14'd 4454: out = 14'h3ADB;
            14'd 4455: out = 14'h3AD8;
            14'd 4456: out = 14'h3AD4;
            14'd 4457: out = 14'h3AD1;
            14'd 4458: out = 14'h3ACE;
            14'd 4459: out = 14'h3ACA;
            14'd 4460: out = 14'h3AC7;
            14'd 4461: out = 14'h3AC3;
            14'd 4462: out = 14'h3AC0;
            14'd 4463: out = 14'h3ABD;
            14'd 4464: out = 14'h3AB9;
            14'd 4465: out = 14'h3AB6;
            14'd 4466: out = 14'h3AB3;
            14'd 4467: out = 14'h3AAF;
            14'd 4468: out = 14'h3AAC;
            14'd 4469: out = 14'h3AA9;
            14'd 4470: out = 14'h3AA5;
            14'd 4471: out = 14'h3AA2;
            14'd 4472: out = 14'h3A9E;
            14'd 4473: out = 14'h3A9B;
            14'd 4474: out = 14'h3A98;
            14'd 4475: out = 14'h3A94;
            14'd 4476: out = 14'h3A91;
            14'd 4477: out = 14'h3A8E;
            14'd 4478: out = 14'h3A8A;
            14'd 4479: out = 14'h3A87;
            14'd 4480: out = 14'h3A84;
            14'd 4481: out = 14'h3A80;
            14'd 4482: out = 14'h3A7D;
            14'd 4483: out = 14'h3A7A;
            14'd 4484: out = 14'h3A76;
            14'd 4485: out = 14'h3A73;
            14'd 4486: out = 14'h3A70;
            14'd 4487: out = 14'h3A6C;
            14'd 4488: out = 14'h3A69;
            14'd 4489: out = 14'h3A66;
            14'd 4490: out = 14'h3A62;
            14'd 4491: out = 14'h3A5F;
            14'd 4492: out = 14'h3A5C;
            14'd 4493: out = 14'h3A58;
            14'd 4494: out = 14'h3A55;
            14'd 4495: out = 14'h3A52;
            14'd 4496: out = 14'h3A4E;
            14'd 4497: out = 14'h3A4B;
            14'd 4498: out = 14'h3A48;
            14'd 4499: out = 14'h3A44;
            14'd 4500: out = 14'h3A41;
            14'd 4501: out = 14'h3A3E;
            14'd 4502: out = 14'h3A3A;
            14'd 4503: out = 14'h3A37;
            14'd 4504: out = 14'h3A34;
            14'd 4505: out = 14'h3A31;
            14'd 4506: out = 14'h3A2D;
            14'd 4507: out = 14'h3A2A;
            14'd 4508: out = 14'h3A27;
            14'd 4509: out = 14'h3A23;
            14'd 4510: out = 14'h3A20;
            14'd 4511: out = 14'h3A1D;
            14'd 4512: out = 14'h3A19;
            14'd 4513: out = 14'h3A16;
            14'd 4514: out = 14'h3A13;
            14'd 4515: out = 14'h3A10;
            14'd 4516: out = 14'h3A0C;
            14'd 4517: out = 14'h3A09;
            14'd 4518: out = 14'h3A06;
            14'd 4519: out = 14'h3A02;
            14'd 4520: out = 14'h39FF;
            14'd 4521: out = 14'h39FC;
            14'd 4522: out = 14'h39F9;
            14'd 4523: out = 14'h39F5;
            14'd 4524: out = 14'h39F2;
            14'd 4525: out = 14'h39EF;
            14'd 4526: out = 14'h39EB;
            14'd 4527: out = 14'h39E8;
            14'd 4528: out = 14'h39E5;
            14'd 4529: out = 14'h39E2;
            14'd 4530: out = 14'h39DE;
            14'd 4531: out = 14'h39DB;
            14'd 4532: out = 14'h39D8;
            14'd 4533: out = 14'h39D5;
            14'd 4534: out = 14'h39D1;
            14'd 4535: out = 14'h39CE;
            14'd 4536: out = 14'h39CB;
            14'd 4537: out = 14'h39C7;
            14'd 4538: out = 14'h39C4;
            14'd 4539: out = 14'h39C1;
            14'd 4540: out = 14'h39BE;
            14'd 4541: out = 14'h39BA;
            14'd 4542: out = 14'h39B7;
            14'd 4543: out = 14'h39B4;
            14'd 4544: out = 14'h39B1;
            14'd 4545: out = 14'h39AD;
            14'd 4546: out = 14'h39AA;
            14'd 4547: out = 14'h39A7;
            14'd 4548: out = 14'h39A4;
            14'd 4549: out = 14'h39A0;
            14'd 4550: out = 14'h399D;
            14'd 4551: out = 14'h399A;
            14'd 4552: out = 14'h3997;
            14'd 4553: out = 14'h3993;
            14'd 4554: out = 14'h3990;
            14'd 4555: out = 14'h398D;
            14'd 4556: out = 14'h398A;
            14'd 4557: out = 14'h3987;
            14'd 4558: out = 14'h3983;
            14'd 4559: out = 14'h3980;
            14'd 4560: out = 14'h397D;
            14'd 4561: out = 14'h397A;
            14'd 4562: out = 14'h3976;
            14'd 4563: out = 14'h3973;
            14'd 4564: out = 14'h3970;
            14'd 4565: out = 14'h396D;
            14'd 4566: out = 14'h396A;
            14'd 4567: out = 14'h3966;
            14'd 4568: out = 14'h3963;
            14'd 4569: out = 14'h3960;
            14'd 4570: out = 14'h395D;
            14'd 4571: out = 14'h3959;
            14'd 4572: out = 14'h3956;
            14'd 4573: out = 14'h3953;
            14'd 4574: out = 14'h3950;
            14'd 4575: out = 14'h394D;
            14'd 4576: out = 14'h3949;
            14'd 4577: out = 14'h3946;
            14'd 4578: out = 14'h3943;
            14'd 4579: out = 14'h3940;
            14'd 4580: out = 14'h393D;
            14'd 4581: out = 14'h3939;
            14'd 4582: out = 14'h3936;
            14'd 4583: out = 14'h3933;
            14'd 4584: out = 14'h3930;
            14'd 4585: out = 14'h392D;
            14'd 4586: out = 14'h3929;
            14'd 4587: out = 14'h3926;
            14'd 4588: out = 14'h3923;
            14'd 4589: out = 14'h3920;
            14'd 4590: out = 14'h391D;
            14'd 4591: out = 14'h3919;
            14'd 4592: out = 14'h3916;
            14'd 4593: out = 14'h3913;
            14'd 4594: out = 14'h3910;
            14'd 4595: out = 14'h390D;
            14'd 4596: out = 14'h390A;
            14'd 4597: out = 14'h3906;
            14'd 4598: out = 14'h3903;
            14'd 4599: out = 14'h3900;
            14'd 4600: out = 14'h38FD;
            14'd 4601: out = 14'h38FA;
            14'd 4602: out = 14'h38F7;
            14'd 4603: out = 14'h38F3;
            14'd 4604: out = 14'h38F0;
            14'd 4605: out = 14'h38ED;
            14'd 4606: out = 14'h38EA;
            14'd 4607: out = 14'h38E7;
            14'd 4608: out = 14'h38E4;
            14'd 4609: out = 14'h38E0;
            14'd 4610: out = 14'h38DD;
            14'd 4611: out = 14'h38DA;
            14'd 4612: out = 14'h38D7;
            14'd 4613: out = 14'h38D4;
            14'd 4614: out = 14'h38D1;
            14'd 4615: out = 14'h38CD;
            14'd 4616: out = 14'h38CA;
            14'd 4617: out = 14'h38C7;
            14'd 4618: out = 14'h38C4;
            14'd 4619: out = 14'h38C1;
            14'd 4620: out = 14'h38BE;
            14'd 4621: out = 14'h38BB;
            14'd 4622: out = 14'h38B7;
            14'd 4623: out = 14'h38B4;
            14'd 4624: out = 14'h38B1;
            14'd 4625: out = 14'h38AE;
            14'd 4626: out = 14'h38AB;
            14'd 4627: out = 14'h38A8;
            14'd 4628: out = 14'h38A5;
            14'd 4629: out = 14'h38A1;
            14'd 4630: out = 14'h389E;
            14'd 4631: out = 14'h389B;
            14'd 4632: out = 14'h3898;
            14'd 4633: out = 14'h3895;
            14'd 4634: out = 14'h3892;
            14'd 4635: out = 14'h388F;
            14'd 4636: out = 14'h388C;
            14'd 4637: out = 14'h3888;
            14'd 4638: out = 14'h3885;
            14'd 4639: out = 14'h3882;
            14'd 4640: out = 14'h387F;
            14'd 4641: out = 14'h387C;
            14'd 4642: out = 14'h3879;
            14'd 4643: out = 14'h3876;
            14'd 4644: out = 14'h3873;
            14'd 4645: out = 14'h3870;
            14'd 4646: out = 14'h386C;
            14'd 4647: out = 14'h3869;
            14'd 4648: out = 14'h3866;
            14'd 4649: out = 14'h3863;
            14'd 4650: out = 14'h3860;
            14'd 4651: out = 14'h385D;
            14'd 4652: out = 14'h385A;
            14'd 4653: out = 14'h3857;
            14'd 4654: out = 14'h3854;
            14'd 4655: out = 14'h3851;
            14'd 4656: out = 14'h384D;
            14'd 4657: out = 14'h384A;
            14'd 4658: out = 14'h3847;
            14'd 4659: out = 14'h3844;
            14'd 4660: out = 14'h3841;
            14'd 4661: out = 14'h383E;
            14'd 4662: out = 14'h383B;
            14'd 4663: out = 14'h3838;
            14'd 4664: out = 14'h3835;
            14'd 4665: out = 14'h3832;
            14'd 4666: out = 14'h382F;
            14'd 4667: out = 14'h382B;
            14'd 4668: out = 14'h3828;
            14'd 4669: out = 14'h3825;
            14'd 4670: out = 14'h3822;
            14'd 4671: out = 14'h381F;
            14'd 4672: out = 14'h381C;
            14'd 4673: out = 14'h3819;
            14'd 4674: out = 14'h3816;
            14'd 4675: out = 14'h3813;
            14'd 4676: out = 14'h3810;
            14'd 4677: out = 14'h380D;
            14'd 4678: out = 14'h380A;
            14'd 4679: out = 14'h3807;
            14'd 4680: out = 14'h3804;
            14'd 4681: out = 14'h3800;
            14'd 4682: out = 14'h37FD;
            14'd 4683: out = 14'h37FA;
            14'd 4684: out = 14'h37F7;
            14'd 4685: out = 14'h37F4;
            14'd 4686: out = 14'h37F1;
            14'd 4687: out = 14'h37EE;
            14'd 4688: out = 14'h37EB;
            14'd 4689: out = 14'h37E8;
            14'd 4690: out = 14'h37E5;
            14'd 4691: out = 14'h37E2;
            14'd 4692: out = 14'h37DF;
            14'd 4693: out = 14'h37DC;
            14'd 4694: out = 14'h37D9;
            14'd 4695: out = 14'h37D6;
            14'd 4696: out = 14'h37D3;
            14'd 4697: out = 14'h37D0;
            14'd 4698: out = 14'h37CD;
            14'd 4699: out = 14'h37CA;
            14'd 4700: out = 14'h37C6;
            14'd 4701: out = 14'h37C3;
            14'd 4702: out = 14'h37C0;
            14'd 4703: out = 14'h37BD;
            14'd 4704: out = 14'h37BA;
            14'd 4705: out = 14'h37B7;
            14'd 4706: out = 14'h37B4;
            14'd 4707: out = 14'h37B1;
            14'd 4708: out = 14'h37AE;
            14'd 4709: out = 14'h37AB;
            14'd 4710: out = 14'h37A8;
            14'd 4711: out = 14'h37A5;
            14'd 4712: out = 14'h37A2;
            14'd 4713: out = 14'h379F;
            14'd 4714: out = 14'h379C;
            14'd 4715: out = 14'h3799;
            14'd 4716: out = 14'h3796;
            14'd 4717: out = 14'h3793;
            14'd 4718: out = 14'h3790;
            14'd 4719: out = 14'h378D;
            14'd 4720: out = 14'h378A;
            14'd 4721: out = 14'h3787;
            14'd 4722: out = 14'h3784;
            14'd 4723: out = 14'h3781;
            14'd 4724: out = 14'h377E;
            14'd 4725: out = 14'h377B;
            14'd 4726: out = 14'h3778;
            14'd 4727: out = 14'h3775;
            14'd 4728: out = 14'h3772;
            14'd 4729: out = 14'h376F;
            14'd 4730: out = 14'h376C;
            14'd 4731: out = 14'h3769;
            14'd 4732: out = 14'h3766;
            14'd 4733: out = 14'h3763;
            14'd 4734: out = 14'h3760;
            14'd 4735: out = 14'h375D;
            14'd 4736: out = 14'h375A;
            14'd 4737: out = 14'h3757;
            14'd 4738: out = 14'h3754;
            14'd 4739: out = 14'h3751;
            14'd 4740: out = 14'h374E;
            14'd 4741: out = 14'h374B;
            14'd 4742: out = 14'h3748;
            14'd 4743: out = 14'h3745;
            14'd 4744: out = 14'h3742;
            14'd 4745: out = 14'h373F;
            14'd 4746: out = 14'h373C;
            14'd 4747: out = 14'h3739;
            14'd 4748: out = 14'h3736;
            14'd 4749: out = 14'h3733;
            14'd 4750: out = 14'h3730;
            14'd 4751: out = 14'h372D;
            14'd 4752: out = 14'h372A;
            14'd 4753: out = 14'h3727;
            14'd 4754: out = 14'h3724;
            14'd 4755: out = 14'h3721;
            14'd 4756: out = 14'h371E;
            14'd 4757: out = 14'h371B;
            14'd 4758: out = 14'h3718;
            14'd 4759: out = 14'h3715;
            14'd 4760: out = 14'h3713;
            14'd 4761: out = 14'h3710;
            14'd 4762: out = 14'h370D;
            14'd 4763: out = 14'h370A;
            14'd 4764: out = 14'h3707;
            14'd 4765: out = 14'h3704;
            14'd 4766: out = 14'h3701;
            14'd 4767: out = 14'h36FE;
            14'd 4768: out = 14'h36FB;
            14'd 4769: out = 14'h36F8;
            14'd 4770: out = 14'h36F5;
            14'd 4771: out = 14'h36F2;
            14'd 4772: out = 14'h36EF;
            14'd 4773: out = 14'h36EC;
            14'd 4774: out = 14'h36E9;
            14'd 4775: out = 14'h36E6;
            14'd 4776: out = 14'h36E3;
            14'd 4777: out = 14'h36E0;
            14'd 4778: out = 14'h36DD;
            14'd 4779: out = 14'h36DA;
            14'd 4780: out = 14'h36D8;
            14'd 4781: out = 14'h36D5;
            14'd 4782: out = 14'h36D2;
            14'd 4783: out = 14'h36CF;
            14'd 4784: out = 14'h36CC;
            14'd 4785: out = 14'h36C9;
            14'd 4786: out = 14'h36C6;
            14'd 4787: out = 14'h36C3;
            14'd 4788: out = 14'h36C0;
            14'd 4789: out = 14'h36BD;
            14'd 4790: out = 14'h36BA;
            14'd 4791: out = 14'h36B7;
            14'd 4792: out = 14'h36B4;
            14'd 4793: out = 14'h36B1;
            14'd 4794: out = 14'h36AF;
            14'd 4795: out = 14'h36AC;
            14'd 4796: out = 14'h36A9;
            14'd 4797: out = 14'h36A6;
            14'd 4798: out = 14'h36A3;
            14'd 4799: out = 14'h36A0;
            14'd 4800: out = 14'h369D;
            14'd 4801: out = 14'h369A;
            14'd 4802: out = 14'h3697;
            14'd 4803: out = 14'h3694;
            14'd 4804: out = 14'h3691;
            14'd 4805: out = 14'h368E;
            14'd 4806: out = 14'h368C;
            14'd 4807: out = 14'h3689;
            14'd 4808: out = 14'h3686;
            14'd 4809: out = 14'h3683;
            14'd 4810: out = 14'h3680;
            14'd 4811: out = 14'h367D;
            14'd 4812: out = 14'h367A;
            14'd 4813: out = 14'h3677;
            14'd 4814: out = 14'h3674;
            14'd 4815: out = 14'h3671;
            14'd 4816: out = 14'h366F;
            14'd 4817: out = 14'h366C;
            14'd 4818: out = 14'h3669;
            14'd 4819: out = 14'h3666;
            14'd 4820: out = 14'h3663;
            14'd 4821: out = 14'h3660;
            14'd 4822: out = 14'h365D;
            14'd 4823: out = 14'h365A;
            14'd 4824: out = 14'h3657;
            14'd 4825: out = 14'h3655;
            14'd 4826: out = 14'h3652;
            14'd 4827: out = 14'h364F;
            14'd 4828: out = 14'h364C;
            14'd 4829: out = 14'h3649;
            14'd 4830: out = 14'h3646;
            14'd 4831: out = 14'h3643;
            14'd 4832: out = 14'h3640;
            14'd 4833: out = 14'h363E;
            14'd 4834: out = 14'h363B;
            14'd 4835: out = 14'h3638;
            14'd 4836: out = 14'h3635;
            14'd 4837: out = 14'h3632;
            14'd 4838: out = 14'h362F;
            14'd 4839: out = 14'h362C;
            14'd 4840: out = 14'h3629;
            14'd 4841: out = 14'h3627;
            14'd 4842: out = 14'h3624;
            14'd 4843: out = 14'h3621;
            14'd 4844: out = 14'h361E;
            14'd 4845: out = 14'h361B;
            14'd 4846: out = 14'h3618;
            14'd 4847: out = 14'h3615;
            14'd 4848: out = 14'h3613;
            14'd 4849: out = 14'h3610;
            14'd 4850: out = 14'h360D;
            14'd 4851: out = 14'h360A;
            14'd 4852: out = 14'h3607;
            14'd 4853: out = 14'h3604;
            14'd 4854: out = 14'h3601;
            14'd 4855: out = 14'h35FF;
            14'd 4856: out = 14'h35FC;
            14'd 4857: out = 14'h35F9;
            14'd 4858: out = 14'h35F6;
            14'd 4859: out = 14'h35F3;
            14'd 4860: out = 14'h35F0;
            14'd 4861: out = 14'h35EE;
            14'd 4862: out = 14'h35EB;
            14'd 4863: out = 14'h35E8;
            14'd 4864: out = 14'h35E5;
            14'd 4865: out = 14'h35E2;
            14'd 4866: out = 14'h35DF;
            14'd 4867: out = 14'h35DD;
            14'd 4868: out = 14'h35DA;
            14'd 4869: out = 14'h35D7;
            14'd 4870: out = 14'h35D4;
            14'd 4871: out = 14'h35D1;
            14'd 4872: out = 14'h35CE;
            14'd 4873: out = 14'h35CC;
            14'd 4874: out = 14'h35C9;
            14'd 4875: out = 14'h35C6;
            14'd 4876: out = 14'h35C3;
            14'd 4877: out = 14'h35C0;
            14'd 4878: out = 14'h35BD;
            14'd 4879: out = 14'h35BB;
            14'd 4880: out = 14'h35B8;
            14'd 4881: out = 14'h35B5;
            14'd 4882: out = 14'h35B2;
            14'd 4883: out = 14'h35AF;
            14'd 4884: out = 14'h35AD;
            14'd 4885: out = 14'h35AA;
            14'd 4886: out = 14'h35A7;
            14'd 4887: out = 14'h35A4;
            14'd 4888: out = 14'h35A1;
            14'd 4889: out = 14'h359F;
            14'd 4890: out = 14'h359C;
            14'd 4891: out = 14'h3599;
            14'd 4892: out = 14'h3596;
            14'd 4893: out = 14'h3593;
            14'd 4894: out = 14'h3590;
            14'd 4895: out = 14'h358E;
            14'd 4896: out = 14'h358B;
            14'd 4897: out = 14'h3588;
            14'd 4898: out = 14'h3585;
            14'd 4899: out = 14'h3582;
            14'd 4900: out = 14'h3580;
            14'd 4901: out = 14'h357D;
            14'd 4902: out = 14'h357A;
            14'd 4903: out = 14'h3577;
            14'd 4904: out = 14'h3575;
            14'd 4905: out = 14'h3572;
            14'd 4906: out = 14'h356F;
            14'd 4907: out = 14'h356C;
            14'd 4908: out = 14'h3569;
            14'd 4909: out = 14'h3567;
            14'd 4910: out = 14'h3564;
            14'd 4911: out = 14'h3561;
            14'd 4912: out = 14'h355E;
            14'd 4913: out = 14'h355B;
            14'd 4914: out = 14'h3559;
            14'd 4915: out = 14'h3556;
            14'd 4916: out = 14'h3553;
            14'd 4917: out = 14'h3550;
            14'd 4918: out = 14'h354E;
            14'd 4919: out = 14'h354B;
            14'd 4920: out = 14'h3548;
            14'd 4921: out = 14'h3545;
            14'd 4922: out = 14'h3542;
            14'd 4923: out = 14'h3540;
            14'd 4924: out = 14'h353D;
            14'd 4925: out = 14'h353A;
            14'd 4926: out = 14'h3537;
            14'd 4927: out = 14'h3535;
            14'd 4928: out = 14'h3532;
            14'd 4929: out = 14'h352F;
            14'd 4930: out = 14'h352C;
            14'd 4931: out = 14'h352A;
            14'd 4932: out = 14'h3527;
            14'd 4933: out = 14'h3524;
            14'd 4934: out = 14'h3521;
            14'd 4935: out = 14'h351F;
            14'd 4936: out = 14'h351C;
            14'd 4937: out = 14'h3519;
            14'd 4938: out = 14'h3516;
            14'd 4939: out = 14'h3514;
            14'd 4940: out = 14'h3511;
            14'd 4941: out = 14'h350E;
            14'd 4942: out = 14'h350B;
            14'd 4943: out = 14'h3509;
            14'd 4944: out = 14'h3506;
            14'd 4945: out = 14'h3503;
            14'd 4946: out = 14'h3500;
            14'd 4947: out = 14'h34FE;
            14'd 4948: out = 14'h34FB;
            14'd 4949: out = 14'h34F8;
            14'd 4950: out = 14'h34F5;
            14'd 4951: out = 14'h34F3;
            14'd 4952: out = 14'h34F0;
            14'd 4953: out = 14'h34ED;
            14'd 4954: out = 14'h34EA;
            14'd 4955: out = 14'h34E8;
            14'd 4956: out = 14'h34E5;
            14'd 4957: out = 14'h34E2;
            14'd 4958: out = 14'h34DF;
            14'd 4959: out = 14'h34DD;
            14'd 4960: out = 14'h34DA;
            14'd 4961: out = 14'h34D7;
            14'd 4962: out = 14'h34D5;
            14'd 4963: out = 14'h34D2;
            14'd 4964: out = 14'h34CF;
            14'd 4965: out = 14'h34CC;
            14'd 4966: out = 14'h34CA;
            14'd 4967: out = 14'h34C7;
            14'd 4968: out = 14'h34C4;
            14'd 4969: out = 14'h34C2;
            14'd 4970: out = 14'h34BF;
            14'd 4971: out = 14'h34BC;
            14'd 4972: out = 14'h34B9;
            14'd 4973: out = 14'h34B7;
            14'd 4974: out = 14'h34B4;
            14'd 4975: out = 14'h34B1;
            14'd 4976: out = 14'h34AF;
            14'd 4977: out = 14'h34AC;
            14'd 4978: out = 14'h34A9;
            14'd 4979: out = 14'h34A6;
            14'd 4980: out = 14'h34A4;
            14'd 4981: out = 14'h34A1;
            14'd 4982: out = 14'h349E;
            14'd 4983: out = 14'h349C;
            14'd 4984: out = 14'h3499;
            14'd 4985: out = 14'h3496;
            14'd 4986: out = 14'h3493;
            14'd 4987: out = 14'h3491;
            14'd 4988: out = 14'h348E;
            14'd 4989: out = 14'h348B;
            14'd 4990: out = 14'h3489;
            14'd 4991: out = 14'h3486;
            14'd 4992: out = 14'h3483;
            14'd 4993: out = 14'h3481;
            14'd 4994: out = 14'h347E;
            14'd 4995: out = 14'h347B;
            14'd 4996: out = 14'h3479;
            14'd 4997: out = 14'h3476;
            14'd 4998: out = 14'h3473;
            14'd 4999: out = 14'h3470;
            14'd 5000: out = 14'h346E;
            14'd 5001: out = 14'h346B;
            14'd 5002: out = 14'h3468;
            14'd 5003: out = 14'h3466;
            14'd 5004: out = 14'h3463;
            14'd 5005: out = 14'h3460;
            14'd 5006: out = 14'h345E;
            14'd 5007: out = 14'h345B;
            14'd 5008: out = 14'h3458;
            14'd 5009: out = 14'h3456;
            14'd 5010: out = 14'h3453;
            14'd 5011: out = 14'h3450;
            14'd 5012: out = 14'h344E;
            14'd 5013: out = 14'h344B;
            14'd 5014: out = 14'h3448;
            14'd 5015: out = 14'h3446;
            14'd 5016: out = 14'h3443;
            14'd 5017: out = 14'h3440;
            14'd 5018: out = 14'h343E;
            14'd 5019: out = 14'h343B;
            14'd 5020: out = 14'h3438;
            14'd 5021: out = 14'h3436;
            14'd 5022: out = 14'h3433;
            14'd 5023: out = 14'h3430;
            14'd 5024: out = 14'h342E;
            14'd 5025: out = 14'h342B;
            14'd 5026: out = 14'h3428;
            14'd 5027: out = 14'h3426;
            14'd 5028: out = 14'h3423;
            14'd 5029: out = 14'h3420;
            14'd 5030: out = 14'h341E;
            14'd 5031: out = 14'h341B;
            14'd 5032: out = 14'h3418;
            14'd 5033: out = 14'h3416;
            14'd 5034: out = 14'h3413;
            14'd 5035: out = 14'h3410;
            14'd 5036: out = 14'h340E;
            14'd 5037: out = 14'h340B;
            14'd 5038: out = 14'h3409;
            14'd 5039: out = 14'h3406;
            14'd 5040: out = 14'h3403;
            14'd 5041: out = 14'h3401;
            14'd 5042: out = 14'h33FE;
            14'd 5043: out = 14'h33FB;
            14'd 5044: out = 14'h33F9;
            14'd 5045: out = 14'h33F6;
            14'd 5046: out = 14'h33F3;
            14'd 5047: out = 14'h33F1;
            14'd 5048: out = 14'h33EE;
            14'd 5049: out = 14'h33EC;
            14'd 5050: out = 14'h33E9;
            14'd 5051: out = 14'h33E6;
            14'd 5052: out = 14'h33E4;
            14'd 5053: out = 14'h33E1;
            14'd 5054: out = 14'h33DE;
            14'd 5055: out = 14'h33DC;
            14'd 5056: out = 14'h33D9;
            14'd 5057: out = 14'h33D6;
            14'd 5058: out = 14'h33D4;
            14'd 5059: out = 14'h33D1;
            14'd 5060: out = 14'h33CF;
            14'd 5061: out = 14'h33CC;
            14'd 5062: out = 14'h33C9;
            14'd 5063: out = 14'h33C7;
            14'd 5064: out = 14'h33C4;
            14'd 5065: out = 14'h33C2;
            14'd 5066: out = 14'h33BF;
            14'd 5067: out = 14'h33BC;
            14'd 5068: out = 14'h33BA;
            14'd 5069: out = 14'h33B7;
            14'd 5070: out = 14'h33B4;
            14'd 5071: out = 14'h33B2;
            14'd 5072: out = 14'h33AF;
            14'd 5073: out = 14'h33AD;
            14'd 5074: out = 14'h33AA;
            14'd 5075: out = 14'h33A7;
            14'd 5076: out = 14'h33A5;
            14'd 5077: out = 14'h33A2;
            14'd 5078: out = 14'h33A0;
            14'd 5079: out = 14'h339D;
            14'd 5080: out = 14'h339A;
            14'd 5081: out = 14'h3398;
            14'd 5082: out = 14'h3395;
            14'd 5083: out = 14'h3393;
            14'd 5084: out = 14'h3390;
            14'd 5085: out = 14'h338D;
            14'd 5086: out = 14'h338B;
            14'd 5087: out = 14'h3388;
            14'd 5088: out = 14'h3386;
            14'd 5089: out = 14'h3383;
            14'd 5090: out = 14'h3380;
            14'd 5091: out = 14'h337E;
            14'd 5092: out = 14'h337B;
            14'd 5093: out = 14'h3379;
            14'd 5094: out = 14'h3376;
            14'd 5095: out = 14'h3374;
            14'd 5096: out = 14'h3371;
            14'd 5097: out = 14'h336E;
            14'd 5098: out = 14'h336C;
            14'd 5099: out = 14'h3369;
            14'd 5100: out = 14'h3367;
            14'd 5101: out = 14'h3364;
            14'd 5102: out = 14'h3361;
            14'd 5103: out = 14'h335F;
            14'd 5104: out = 14'h335C;
            14'd 5105: out = 14'h335A;
            14'd 5106: out = 14'h3357;
            14'd 5107: out = 14'h3355;
            14'd 5108: out = 14'h3352;
            14'd 5109: out = 14'h334F;
            14'd 5110: out = 14'h334D;
            14'd 5111: out = 14'h334A;
            14'd 5112: out = 14'h3348;
            14'd 5113: out = 14'h3345;
            14'd 5114: out = 14'h3343;
            14'd 5115: out = 14'h3340;
            14'd 5116: out = 14'h333D;
            14'd 5117: out = 14'h333B;
            14'd 5118: out = 14'h3338;
            14'd 5119: out = 14'h3336;
            14'd 5120: out = 14'h3333;
            14'd 5121: out = 14'h3331;
            14'd 5122: out = 14'h332E;
            14'd 5123: out = 14'h332C;
            14'd 5124: out = 14'h3329;
            14'd 5125: out = 14'h3326;
            14'd 5126: out = 14'h3324;
            14'd 5127: out = 14'h3321;
            14'd 5128: out = 14'h331F;
            14'd 5129: out = 14'h331C;
            14'd 5130: out = 14'h331A;
            14'd 5131: out = 14'h3317;
            14'd 5132: out = 14'h3315;
            14'd 5133: out = 14'h3312;
            14'd 5134: out = 14'h330F;
            14'd 5135: out = 14'h330D;
            14'd 5136: out = 14'h330A;
            14'd 5137: out = 14'h3308;
            14'd 5138: out = 14'h3305;
            14'd 5139: out = 14'h3303;
            14'd 5140: out = 14'h3300;
            14'd 5141: out = 14'h32FE;
            14'd 5142: out = 14'h32FB;
            14'd 5143: out = 14'h32F9;
            14'd 5144: out = 14'h32F6;
            14'd 5145: out = 14'h32F4;
            14'd 5146: out = 14'h32F1;
            14'd 5147: out = 14'h32EE;
            14'd 5148: out = 14'h32EC;
            14'd 5149: out = 14'h32E9;
            14'd 5150: out = 14'h32E7;
            14'd 5151: out = 14'h32E4;
            14'd 5152: out = 14'h32E2;
            14'd 5153: out = 14'h32DF;
            14'd 5154: out = 14'h32DD;
            14'd 5155: out = 14'h32DA;
            14'd 5156: out = 14'h32D8;
            14'd 5157: out = 14'h32D5;
            14'd 5158: out = 14'h32D3;
            14'd 5159: out = 14'h32D0;
            14'd 5160: out = 14'h32CE;
            14'd 5161: out = 14'h32CB;
            14'd 5162: out = 14'h32C9;
            14'd 5163: out = 14'h32C6;
            14'd 5164: out = 14'h32C4;
            14'd 5165: out = 14'h32C1;
            14'd 5166: out = 14'h32BE;
            14'd 5167: out = 14'h32BC;
            14'd 5168: out = 14'h32B9;
            14'd 5169: out = 14'h32B7;
            14'd 5170: out = 14'h32B4;
            14'd 5171: out = 14'h32B2;
            14'd 5172: out = 14'h32AF;
            14'd 5173: out = 14'h32AD;
            14'd 5174: out = 14'h32AA;
            14'd 5175: out = 14'h32A8;
            14'd 5176: out = 14'h32A5;
            14'd 5177: out = 14'h32A3;
            14'd 5178: out = 14'h32A0;
            14'd 5179: out = 14'h329E;
            14'd 5180: out = 14'h329B;
            14'd 5181: out = 14'h3299;
            14'd 5182: out = 14'h3296;
            14'd 5183: out = 14'h3294;
            14'd 5184: out = 14'h3291;
            14'd 5185: out = 14'h328F;
            14'd 5186: out = 14'h328C;
            14'd 5187: out = 14'h328A;
            14'd 5188: out = 14'h3287;
            14'd 5189: out = 14'h3285;
            14'd 5190: out = 14'h3282;
            14'd 5191: out = 14'h3280;
            14'd 5192: out = 14'h327D;
            14'd 5193: out = 14'h327B;
            14'd 5194: out = 14'h3278;
            14'd 5195: out = 14'h3276;
            14'd 5196: out = 14'h3273;
            14'd 5197: out = 14'h3271;
            14'd 5198: out = 14'h326F;
            14'd 5199: out = 14'h326C;
            14'd 5200: out = 14'h326A;
            14'd 5201: out = 14'h3267;
            14'd 5202: out = 14'h3265;
            14'd 5203: out = 14'h3262;
            14'd 5204: out = 14'h3260;
            14'd 5205: out = 14'h325D;
            14'd 5206: out = 14'h325B;
            14'd 5207: out = 14'h3258;
            14'd 5208: out = 14'h3256;
            14'd 5209: out = 14'h3253;
            14'd 5210: out = 14'h3251;
            14'd 5211: out = 14'h324E;
            14'd 5212: out = 14'h324C;
            14'd 5213: out = 14'h3249;
            14'd 5214: out = 14'h3247;
            14'd 5215: out = 14'h3244;
            14'd 5216: out = 14'h3242;
            14'd 5217: out = 14'h323F;
            14'd 5218: out = 14'h323D;
            14'd 5219: out = 14'h323B;
            14'd 5220: out = 14'h3238;
            14'd 5221: out = 14'h3236;
            14'd 5222: out = 14'h3233;
            14'd 5223: out = 14'h3231;
            14'd 5224: out = 14'h322E;
            14'd 5225: out = 14'h322C;
            14'd 5226: out = 14'h3229;
            14'd 5227: out = 14'h3227;
            14'd 5228: out = 14'h3224;
            14'd 5229: out = 14'h3222;
            14'd 5230: out = 14'h3220;
            14'd 5231: out = 14'h321D;
            14'd 5232: out = 14'h321B;
            14'd 5233: out = 14'h3218;
            14'd 5234: out = 14'h3216;
            14'd 5235: out = 14'h3213;
            14'd 5236: out = 14'h3211;
            14'd 5237: out = 14'h320E;
            14'd 5238: out = 14'h320C;
            14'd 5239: out = 14'h3209;
            14'd 5240: out = 14'h3207;
            14'd 5241: out = 14'h3205;
            14'd 5242: out = 14'h3202;
            14'd 5243: out = 14'h3200;
            14'd 5244: out = 14'h31FD;
            14'd 5245: out = 14'h31FB;
            14'd 5246: out = 14'h31F8;
            14'd 5247: out = 14'h31F6;
            14'd 5248: out = 14'h31F4;
            14'd 5249: out = 14'h31F1;
            14'd 5250: out = 14'h31EF;
            14'd 5251: out = 14'h31EC;
            14'd 5252: out = 14'h31EA;
            14'd 5253: out = 14'h31E7;
            14'd 5254: out = 14'h31E5;
            14'd 5255: out = 14'h31E2;
            14'd 5256: out = 14'h31E0;
            14'd 5257: out = 14'h31DE;
            14'd 5258: out = 14'h31DB;
            14'd 5259: out = 14'h31D9;
            14'd 5260: out = 14'h31D6;
            14'd 5261: out = 14'h31D4;
            14'd 5262: out = 14'h31D1;
            14'd 5263: out = 14'h31CF;
            14'd 5264: out = 14'h31CD;
            14'd 5265: out = 14'h31CA;
            14'd 5266: out = 14'h31C8;
            14'd 5267: out = 14'h31C5;
            14'd 5268: out = 14'h31C3;
            14'd 5269: out = 14'h31C1;
            14'd 5270: out = 14'h31BE;
            14'd 5271: out = 14'h31BC;
            14'd 5272: out = 14'h31B9;
            14'd 5273: out = 14'h31B7;
            14'd 5274: out = 14'h31B4;
            14'd 5275: out = 14'h31B2;
            14'd 5276: out = 14'h31B0;
            14'd 5277: out = 14'h31AD;
            14'd 5278: out = 14'h31AB;
            14'd 5279: out = 14'h31A8;
            14'd 5280: out = 14'h31A6;
            14'd 5281: out = 14'h31A4;
            14'd 5282: out = 14'h31A1;
            14'd 5283: out = 14'h319F;
            14'd 5284: out = 14'h319C;
            14'd 5285: out = 14'h319A;
            14'd 5286: out = 14'h3198;
            14'd 5287: out = 14'h3195;
            14'd 5288: out = 14'h3193;
            14'd 5289: out = 14'h3190;
            14'd 5290: out = 14'h318E;
            14'd 5291: out = 14'h318C;
            14'd 5292: out = 14'h3189;
            14'd 5293: out = 14'h3187;
            14'd 5294: out = 14'h3184;
            14'd 5295: out = 14'h3182;
            14'd 5296: out = 14'h3180;
            14'd 5297: out = 14'h317D;
            14'd 5298: out = 14'h317B;
            14'd 5299: out = 14'h3178;
            14'd 5300: out = 14'h3176;
            14'd 5301: out = 14'h3174;
            14'd 5302: out = 14'h3171;
            14'd 5303: out = 14'h316F;
            14'd 5304: out = 14'h316D;
            14'd 5305: out = 14'h316A;
            14'd 5306: out = 14'h3168;
            14'd 5307: out = 14'h3165;
            14'd 5308: out = 14'h3163;
            14'd 5309: out = 14'h3161;
            14'd 5310: out = 14'h315E;
            14'd 5311: out = 14'h315C;
            14'd 5312: out = 14'h3159;
            14'd 5313: out = 14'h3157;
            14'd 5314: out = 14'h3155;
            14'd 5315: out = 14'h3152;
            14'd 5316: out = 14'h3150;
            14'd 5317: out = 14'h314E;
            14'd 5318: out = 14'h314B;
            14'd 5319: out = 14'h3149;
            14'd 5320: out = 14'h3146;
            14'd 5321: out = 14'h3144;
            14'd 5322: out = 14'h3142;
            14'd 5323: out = 14'h313F;
            14'd 5324: out = 14'h313D;
            14'd 5325: out = 14'h313B;
            14'd 5326: out = 14'h3138;
            14'd 5327: out = 14'h3136;
            14'd 5328: out = 14'h3134;
            14'd 5329: out = 14'h3131;
            14'd 5330: out = 14'h312F;
            14'd 5331: out = 14'h312C;
            14'd 5332: out = 14'h312A;
            14'd 5333: out = 14'h3128;
            14'd 5334: out = 14'h3125;
            14'd 5335: out = 14'h3123;
            14'd 5336: out = 14'h3121;
            14'd 5337: out = 14'h311E;
            14'd 5338: out = 14'h311C;
            14'd 5339: out = 14'h311A;
            14'd 5340: out = 14'h3117;
            14'd 5341: out = 14'h3115;
            14'd 5342: out = 14'h3112;
            14'd 5343: out = 14'h3110;
            14'd 5344: out = 14'h310E;
            14'd 5345: out = 14'h310B;
            14'd 5346: out = 14'h3109;
            14'd 5347: out = 14'h3107;
            14'd 5348: out = 14'h3104;
            14'd 5349: out = 14'h3102;
            14'd 5350: out = 14'h3100;
            14'd 5351: out = 14'h30FD;
            14'd 5352: out = 14'h30FB;
            14'd 5353: out = 14'h30F9;
            14'd 5354: out = 14'h30F6;
            14'd 5355: out = 14'h30F4;
            14'd 5356: out = 14'h30F2;
            14'd 5357: out = 14'h30EF;
            14'd 5358: out = 14'h30ED;
            14'd 5359: out = 14'h30EB;
            14'd 5360: out = 14'h30E8;
            14'd 5361: out = 14'h30E6;
            14'd 5362: out = 14'h30E4;
            14'd 5363: out = 14'h30E1;
            14'd 5364: out = 14'h30DF;
            14'd 5365: out = 14'h30DD;
            14'd 5366: out = 14'h30DA;
            14'd 5367: out = 14'h30D8;
            14'd 5368: out = 14'h30D6;
            14'd 5369: out = 14'h30D3;
            14'd 5370: out = 14'h30D1;
            14'd 5371: out = 14'h30CF;
            14'd 5372: out = 14'h30CC;
            14'd 5373: out = 14'h30CA;
            14'd 5374: out = 14'h30C8;
            14'd 5375: out = 14'h30C5;
            14'd 5376: out = 14'h30C3;
            14'd 5377: out = 14'h30C1;
            14'd 5378: out = 14'h30BE;
            14'd 5379: out = 14'h30BC;
            14'd 5380: out = 14'h30BA;
            14'd 5381: out = 14'h30B7;
            14'd 5382: out = 14'h30B5;
            14'd 5383: out = 14'h30B3;
            14'd 5384: out = 14'h30B0;
            14'd 5385: out = 14'h30AE;
            14'd 5386: out = 14'h30AC;
            14'd 5387: out = 14'h30AA;
            14'd 5388: out = 14'h30A7;
            14'd 5389: out = 14'h30A5;
            14'd 5390: out = 14'h30A3;
            14'd 5391: out = 14'h30A0;
            14'd 5392: out = 14'h309E;
            14'd 5393: out = 14'h309C;
            14'd 5394: out = 14'h3099;
            14'd 5395: out = 14'h3097;
            14'd 5396: out = 14'h3095;
            14'd 5397: out = 14'h3092;
            14'd 5398: out = 14'h3090;
            14'd 5399: out = 14'h308E;
            14'd 5400: out = 14'h308C;
            14'd 5401: out = 14'h3089;
            14'd 5402: out = 14'h3087;
            14'd 5403: out = 14'h3085;
            14'd 5404: out = 14'h3082;
            14'd 5405: out = 14'h3080;
            14'd 5406: out = 14'h307E;
            14'd 5407: out = 14'h307B;
            14'd 5408: out = 14'h3079;
            14'd 5409: out = 14'h3077;
            14'd 5410: out = 14'h3075;
            14'd 5411: out = 14'h3072;
            14'd 5412: out = 14'h3070;
            14'd 5413: out = 14'h306E;
            14'd 5414: out = 14'h306B;
            14'd 5415: out = 14'h3069;
            14'd 5416: out = 14'h3067;
            14'd 5417: out = 14'h3065;
            14'd 5418: out = 14'h3062;
            14'd 5419: out = 14'h3060;
            14'd 5420: out = 14'h305E;
            14'd 5421: out = 14'h305B;
            14'd 5422: out = 14'h3059;
            14'd 5423: out = 14'h3057;
            14'd 5424: out = 14'h3055;
            14'd 5425: out = 14'h3052;
            14'd 5426: out = 14'h3050;
            14'd 5427: out = 14'h304E;
            14'd 5428: out = 14'h304B;
            14'd 5429: out = 14'h3049;
            14'd 5430: out = 14'h3047;
            14'd 5431: out = 14'h3045;
            14'd 5432: out = 14'h3042;
            14'd 5433: out = 14'h3040;
            14'd 5434: out = 14'h303E;
            14'd 5435: out = 14'h303C;
            14'd 5436: out = 14'h3039;
            14'd 5437: out = 14'h3037;
            14'd 5438: out = 14'h3035;
            14'd 5439: out = 14'h3032;
            14'd 5440: out = 14'h3030;
            14'd 5441: out = 14'h302E;
            14'd 5442: out = 14'h302C;
            14'd 5443: out = 14'h3029;
            14'd 5444: out = 14'h3027;
            14'd 5445: out = 14'h3025;
            14'd 5446: out = 14'h3023;
            14'd 5447: out = 14'h3020;
            14'd 5448: out = 14'h301E;
            14'd 5449: out = 14'h301C;
            14'd 5450: out = 14'h301A;
            14'd 5451: out = 14'h3017;
            14'd 5452: out = 14'h3015;
            14'd 5453: out = 14'h3013;
            14'd 5454: out = 14'h3011;
            14'd 5455: out = 14'h300E;
            14'd 5456: out = 14'h300C;
            14'd 5457: out = 14'h300A;
            14'd 5458: out = 14'h3008;
            14'd 5459: out = 14'h3005;
            14'd 5460: out = 14'h3003;
            14'd 5461: out = 14'h3001;
            14'd 5462: out = 14'h2FFF;
            14'd 5463: out = 14'h2FFC;
            14'd 5464: out = 14'h2FFA;
            14'd 5465: out = 14'h2FF8;
            14'd 5466: out = 14'h2FF6;
            14'd 5467: out = 14'h2FF3;
            14'd 5468: out = 14'h2FF1;
            14'd 5469: out = 14'h2FEF;
            14'd 5470: out = 14'h2FED;
            14'd 5471: out = 14'h2FEA;
            14'd 5472: out = 14'h2FE8;
            14'd 5473: out = 14'h2FE6;
            14'd 5474: out = 14'h2FE4;
            14'd 5475: out = 14'h2FE1;
            14'd 5476: out = 14'h2FDF;
            14'd 5477: out = 14'h2FDD;
            14'd 5478: out = 14'h2FDB;
            14'd 5479: out = 14'h2FD8;
            14'd 5480: out = 14'h2FD6;
            14'd 5481: out = 14'h2FD4;
            14'd 5482: out = 14'h2FD2;
            14'd 5483: out = 14'h2FCF;
            14'd 5484: out = 14'h2FCD;
            14'd 5485: out = 14'h2FCB;
            14'd 5486: out = 14'h2FC9;
            14'd 5487: out = 14'h2FC7;
            14'd 5488: out = 14'h2FC4;
            14'd 5489: out = 14'h2FC2;
            14'd 5490: out = 14'h2FC0;
            14'd 5491: out = 14'h2FBE;
            14'd 5492: out = 14'h2FBB;
            14'd 5493: out = 14'h2FB9;
            14'd 5494: out = 14'h2FB7;
            14'd 5495: out = 14'h2FB5;
            14'd 5496: out = 14'h2FB2;
            14'd 5497: out = 14'h2FB0;
            14'd 5498: out = 14'h2FAE;
            14'd 5499: out = 14'h2FAC;
            14'd 5500: out = 14'h2FAA;
            14'd 5501: out = 14'h2FA7;
            14'd 5502: out = 14'h2FA5;
            14'd 5503: out = 14'h2FA3;
            14'd 5504: out = 14'h2FA1;
            14'd 5505: out = 14'h2F9F;
            14'd 5506: out = 14'h2F9C;
            14'd 5507: out = 14'h2F9A;
            14'd 5508: out = 14'h2F98;
            14'd 5509: out = 14'h2F96;
            14'd 5510: out = 14'h2F93;
            14'd 5511: out = 14'h2F91;
            14'd 5512: out = 14'h2F8F;
            14'd 5513: out = 14'h2F8D;
            14'd 5514: out = 14'h2F8B;
            14'd 5515: out = 14'h2F88;
            14'd 5516: out = 14'h2F86;
            14'd 5517: out = 14'h2F84;
            14'd 5518: out = 14'h2F82;
            14'd 5519: out = 14'h2F80;
            14'd 5520: out = 14'h2F7D;
            14'd 5521: out = 14'h2F7B;
            14'd 5522: out = 14'h2F79;
            14'd 5523: out = 14'h2F77;
            14'd 5524: out = 14'h2F75;
            14'd 5525: out = 14'h2F72;
            14'd 5526: out = 14'h2F70;
            14'd 5527: out = 14'h2F6E;
            14'd 5528: out = 14'h2F6C;
            14'd 5529: out = 14'h2F6A;
            14'd 5530: out = 14'h2F67;
            14'd 5531: out = 14'h2F65;
            14'd 5532: out = 14'h2F63;
            14'd 5533: out = 14'h2F61;
            14'd 5534: out = 14'h2F5F;
            14'd 5535: out = 14'h2F5C;
            14'd 5536: out = 14'h2F5A;
            14'd 5537: out = 14'h2F58;
            14'd 5538: out = 14'h2F56;
            14'd 5539: out = 14'h2F54;
            14'd 5540: out = 14'h2F52;
            14'd 5541: out = 14'h2F4F;
            14'd 5542: out = 14'h2F4D;
            14'd 5543: out = 14'h2F4B;
            14'd 5544: out = 14'h2F49;
            14'd 5545: out = 14'h2F47;
            14'd 5546: out = 14'h2F44;
            14'd 5547: out = 14'h2F42;
            14'd 5548: out = 14'h2F40;
            14'd 5549: out = 14'h2F3E;
            14'd 5550: out = 14'h2F3C;
            14'd 5551: out = 14'h2F3A;
            14'd 5552: out = 14'h2F37;
            14'd 5553: out = 14'h2F35;
            14'd 5554: out = 14'h2F33;
            14'd 5555: out = 14'h2F31;
            14'd 5556: out = 14'h2F2F;
            14'd 5557: out = 14'h2F2C;
            14'd 5558: out = 14'h2F2A;
            14'd 5559: out = 14'h2F28;
            14'd 5560: out = 14'h2F26;
            14'd 5561: out = 14'h2F24;
            14'd 5562: out = 14'h2F22;
            14'd 5563: out = 14'h2F1F;
            14'd 5564: out = 14'h2F1D;
            14'd 5565: out = 14'h2F1B;
            14'd 5566: out = 14'h2F19;
            14'd 5567: out = 14'h2F17;
            14'd 5568: out = 14'h2F15;
            14'd 5569: out = 14'h2F12;
            14'd 5570: out = 14'h2F10;
            14'd 5571: out = 14'h2F0E;
            14'd 5572: out = 14'h2F0C;
            14'd 5573: out = 14'h2F0A;
            14'd 5574: out = 14'h2F08;
            14'd 5575: out = 14'h2F05;
            14'd 5576: out = 14'h2F03;
            14'd 5577: out = 14'h2F01;
            14'd 5578: out = 14'h2EFF;
            14'd 5579: out = 14'h2EFD;
            14'd 5580: out = 14'h2EFB;
            14'd 5581: out = 14'h2EF9;
            14'd 5582: out = 14'h2EF6;
            14'd 5583: out = 14'h2EF4;
            14'd 5584: out = 14'h2EF2;
            14'd 5585: out = 14'h2EF0;
            14'd 5586: out = 14'h2EEE;
            14'd 5587: out = 14'h2EEC;
            14'd 5588: out = 14'h2EE9;
            14'd 5589: out = 14'h2EE7;
            14'd 5590: out = 14'h2EE5;
            14'd 5591: out = 14'h2EE3;
            14'd 5592: out = 14'h2EE1;
            14'd 5593: out = 14'h2EDF;
            14'd 5594: out = 14'h2EDD;
            14'd 5595: out = 14'h2EDA;
            14'd 5596: out = 14'h2ED8;
            14'd 5597: out = 14'h2ED6;
            14'd 5598: out = 14'h2ED4;
            14'd 5599: out = 14'h2ED2;
            14'd 5600: out = 14'h2ED0;
            14'd 5601: out = 14'h2ECE;
            14'd 5602: out = 14'h2ECB;
            14'd 5603: out = 14'h2EC9;
            14'd 5604: out = 14'h2EC7;
            14'd 5605: out = 14'h2EC5;
            14'd 5606: out = 14'h2EC3;
            14'd 5607: out = 14'h2EC1;
            14'd 5608: out = 14'h2EBF;
            14'd 5609: out = 14'h2EBC;
            14'd 5610: out = 14'h2EBA;
            14'd 5611: out = 14'h2EB8;
            14'd 5612: out = 14'h2EB6;
            14'd 5613: out = 14'h2EB4;
            14'd 5614: out = 14'h2EB2;
            14'd 5615: out = 14'h2EB0;
            14'd 5616: out = 14'h2EAE;
            14'd 5617: out = 14'h2EAB;
            14'd 5618: out = 14'h2EA9;
            14'd 5619: out = 14'h2EA7;
            14'd 5620: out = 14'h2EA5;
            14'd 5621: out = 14'h2EA3;
            14'd 5622: out = 14'h2EA1;
            14'd 5623: out = 14'h2E9F;
            14'd 5624: out = 14'h2E9D;
            14'd 5625: out = 14'h2E9A;
            14'd 5626: out = 14'h2E98;
            14'd 5627: out = 14'h2E96;
            14'd 5628: out = 14'h2E94;
            14'd 5629: out = 14'h2E92;
            14'd 5630: out = 14'h2E90;
            14'd 5631: out = 14'h2E8E;
            14'd 5632: out = 14'h2E8C;
            14'd 5633: out = 14'h2E8A;
            14'd 5634: out = 14'h2E87;
            14'd 5635: out = 14'h2E85;
            14'd 5636: out = 14'h2E83;
            14'd 5637: out = 14'h2E81;
            14'd 5638: out = 14'h2E7F;
            14'd 5639: out = 14'h2E7D;
            14'd 5640: out = 14'h2E7B;
            14'd 5641: out = 14'h2E79;
            14'd 5642: out = 14'h2E77;
            14'd 5643: out = 14'h2E74;
            14'd 5644: out = 14'h2E72;
            14'd 5645: out = 14'h2E70;
            14'd 5646: out = 14'h2E6E;
            14'd 5647: out = 14'h2E6C;
            14'd 5648: out = 14'h2E6A;
            14'd 5649: out = 14'h2E68;
            14'd 5650: out = 14'h2E66;
            14'd 5651: out = 14'h2E64;
            14'd 5652: out = 14'h2E61;
            14'd 5653: out = 14'h2E5F;
            14'd 5654: out = 14'h2E5D;
            14'd 5655: out = 14'h2E5B;
            14'd 5656: out = 14'h2E59;
            14'd 5657: out = 14'h2E57;
            14'd 5658: out = 14'h2E55;
            14'd 5659: out = 14'h2E53;
            14'd 5660: out = 14'h2E51;
            14'd 5661: out = 14'h2E4F;
            14'd 5662: out = 14'h2E4D;
            14'd 5663: out = 14'h2E4A;
            14'd 5664: out = 14'h2E48;
            14'd 5665: out = 14'h2E46;
            14'd 5666: out = 14'h2E44;
            14'd 5667: out = 14'h2E42;
            14'd 5668: out = 14'h2E40;
            14'd 5669: out = 14'h2E3E;
            14'd 5670: out = 14'h2E3C;
            14'd 5671: out = 14'h2E3A;
            14'd 5672: out = 14'h2E38;
            14'd 5673: out = 14'h2E36;
            14'd 5674: out = 14'h2E33;
            14'd 5675: out = 14'h2E31;
            14'd 5676: out = 14'h2E2F;
            14'd 5677: out = 14'h2E2D;
            14'd 5678: out = 14'h2E2B;
            14'd 5679: out = 14'h2E29;
            14'd 5680: out = 14'h2E27;
            14'd 5681: out = 14'h2E25;
            14'd 5682: out = 14'h2E23;
            14'd 5683: out = 14'h2E21;
            14'd 5684: out = 14'h2E1F;
            14'd 5685: out = 14'h2E1D;
            14'd 5686: out = 14'h2E1A;
            14'd 5687: out = 14'h2E18;
            14'd 5688: out = 14'h2E16;
            14'd 5689: out = 14'h2E14;
            14'd 5690: out = 14'h2E12;
            14'd 5691: out = 14'h2E10;
            14'd 5692: out = 14'h2E0E;
            14'd 5693: out = 14'h2E0C;
            14'd 5694: out = 14'h2E0A;
            14'd 5695: out = 14'h2E08;
            14'd 5696: out = 14'h2E06;
            14'd 5697: out = 14'h2E04;
            14'd 5698: out = 14'h2E02;
            14'd 5699: out = 14'h2E00;
            14'd 5700: out = 14'h2DFD;
            14'd 5701: out = 14'h2DFB;
            14'd 5702: out = 14'h2DF9;
            14'd 5703: out = 14'h2DF7;
            14'd 5704: out = 14'h2DF5;
            14'd 5705: out = 14'h2DF3;
            14'd 5706: out = 14'h2DF1;
            14'd 5707: out = 14'h2DEF;
            14'd 5708: out = 14'h2DED;
            14'd 5709: out = 14'h2DEB;
            14'd 5710: out = 14'h2DE9;
            14'd 5711: out = 14'h2DE7;
            14'd 5712: out = 14'h2DE5;
            14'd 5713: out = 14'h2DE3;
            14'd 5714: out = 14'h2DE1;
            14'd 5715: out = 14'h2DDF;
            14'd 5716: out = 14'h2DDD;
            14'd 5717: out = 14'h2DDA;
            14'd 5718: out = 14'h2DD8;
            14'd 5719: out = 14'h2DD6;
            14'd 5720: out = 14'h2DD4;
            14'd 5721: out = 14'h2DD2;
            14'd 5722: out = 14'h2DD0;
            14'd 5723: out = 14'h2DCE;
            14'd 5724: out = 14'h2DCC;
            14'd 5725: out = 14'h2DCA;
            14'd 5726: out = 14'h2DC8;
            14'd 5727: out = 14'h2DC6;
            14'd 5728: out = 14'h2DC4;
            14'd 5729: out = 14'h2DC2;
            14'd 5730: out = 14'h2DC0;
            14'd 5731: out = 14'h2DBE;
            14'd 5732: out = 14'h2DBC;
            14'd 5733: out = 14'h2DBA;
            14'd 5734: out = 14'h2DB8;
            14'd 5735: out = 14'h2DB6;
            14'd 5736: out = 14'h2DB4;
            14'd 5737: out = 14'h2DB2;
            14'd 5738: out = 14'h2DB0;
            14'd 5739: out = 14'h2DAD;
            14'd 5740: out = 14'h2DAB;
            14'd 5741: out = 14'h2DA9;
            14'd 5742: out = 14'h2DA7;
            14'd 5743: out = 14'h2DA5;
            14'd 5744: out = 14'h2DA3;
            14'd 5745: out = 14'h2DA1;
            14'd 5746: out = 14'h2D9F;
            14'd 5747: out = 14'h2D9D;
            14'd 5748: out = 14'h2D9B;
            14'd 5749: out = 14'h2D99;
            14'd 5750: out = 14'h2D97;
            14'd 5751: out = 14'h2D95;
            14'd 5752: out = 14'h2D93;
            14'd 5753: out = 14'h2D91;
            14'd 5754: out = 14'h2D8F;
            14'd 5755: out = 14'h2D8D;
            14'd 5756: out = 14'h2D8B;
            14'd 5757: out = 14'h2D89;
            14'd 5758: out = 14'h2D87;
            14'd 5759: out = 14'h2D85;
            14'd 5760: out = 14'h2D83;
            14'd 5761: out = 14'h2D81;
            14'd 5762: out = 14'h2D7F;
            14'd 5763: out = 14'h2D7D;
            14'd 5764: out = 14'h2D7B;
            14'd 5765: out = 14'h2D79;
            14'd 5766: out = 14'h2D77;
            14'd 5767: out = 14'h2D75;
            14'd 5768: out = 14'h2D73;
            14'd 5769: out = 14'h2D71;
            14'd 5770: out = 14'h2D6F;
            14'd 5771: out = 14'h2D6D;
            14'd 5772: out = 14'h2D6B;
            14'd 5773: out = 14'h2D69;
            14'd 5774: out = 14'h2D67;
            14'd 5775: out = 14'h2D65;
            14'd 5776: out = 14'h2D63;
            14'd 5777: out = 14'h2D61;
            14'd 5778: out = 14'h2D5F;
            14'd 5779: out = 14'h2D5D;
            14'd 5780: out = 14'h2D5B;
            14'd 5781: out = 14'h2D59;
            14'd 5782: out = 14'h2D57;
            14'd 5783: out = 14'h2D55;
            14'd 5784: out = 14'h2D53;
            14'd 5785: out = 14'h2D50;
            14'd 5786: out = 14'h2D4E;
            14'd 5787: out = 14'h2D4C;
            14'd 5788: out = 14'h2D4A;
            14'd 5789: out = 14'h2D48;
            14'd 5790: out = 14'h2D46;
            14'd 5791: out = 14'h2D44;
            14'd 5792: out = 14'h2D42;
            14'd 5793: out = 14'h2D40;
            14'd 5794: out = 14'h2D3E;
            14'd 5795: out = 14'h2D3C;
            14'd 5796: out = 14'h2D3A;
            14'd 5797: out = 14'h2D38;
            14'd 5798: out = 14'h2D36;
            14'd 5799: out = 14'h2D34;
            14'd 5800: out = 14'h2D32;
            14'd 5801: out = 14'h2D30;
            14'd 5802: out = 14'h2D2F;
            14'd 5803: out = 14'h2D2D;
            14'd 5804: out = 14'h2D2B;
            14'd 5805: out = 14'h2D29;
            14'd 5806: out = 14'h2D27;
            14'd 5807: out = 14'h2D25;
            14'd 5808: out = 14'h2D23;
            14'd 5809: out = 14'h2D21;
            14'd 5810: out = 14'h2D1F;
            14'd 5811: out = 14'h2D1D;
            14'd 5812: out = 14'h2D1B;
            14'd 5813: out = 14'h2D19;
            14'd 5814: out = 14'h2D17;
            14'd 5815: out = 14'h2D15;
            14'd 5816: out = 14'h2D13;
            14'd 5817: out = 14'h2D11;
            14'd 5818: out = 14'h2D0F;
            14'd 5819: out = 14'h2D0D;
            14'd 5820: out = 14'h2D0B;
            14'd 5821: out = 14'h2D09;
            14'd 5822: out = 14'h2D07;
            14'd 5823: out = 14'h2D05;
            14'd 5824: out = 14'h2D03;
            14'd 5825: out = 14'h2D01;
            14'd 5826: out = 14'h2CFF;
            14'd 5827: out = 14'h2CFD;
            14'd 5828: out = 14'h2CFB;
            14'd 5829: out = 14'h2CF9;
            14'd 5830: out = 14'h2CF7;
            14'd 5831: out = 14'h2CF5;
            14'd 5832: out = 14'h2CF3;
            14'd 5833: out = 14'h2CF1;
            14'd 5834: out = 14'h2CEF;
            14'd 5835: out = 14'h2CED;
            14'd 5836: out = 14'h2CEB;
            14'd 5837: out = 14'h2CE9;
            14'd 5838: out = 14'h2CE7;
            14'd 5839: out = 14'h2CE5;
            14'd 5840: out = 14'h2CE3;
            14'd 5841: out = 14'h2CE1;
            14'd 5842: out = 14'h2CDF;
            14'd 5843: out = 14'h2CDD;
            14'd 5844: out = 14'h2CDB;
            14'd 5845: out = 14'h2CD9;
            14'd 5846: out = 14'h2CD7;
            14'd 5847: out = 14'h2CD5;
            14'd 5848: out = 14'h2CD4;
            14'd 5849: out = 14'h2CD2;
            14'd 5850: out = 14'h2CD0;
            14'd 5851: out = 14'h2CCE;
            14'd 5852: out = 14'h2CCC;
            14'd 5853: out = 14'h2CCA;
            14'd 5854: out = 14'h2CC8;
            14'd 5855: out = 14'h2CC6;
            14'd 5856: out = 14'h2CC4;
            14'd 5857: out = 14'h2CC2;
            14'd 5858: out = 14'h2CC0;
            14'd 5859: out = 14'h2CBE;
            14'd 5860: out = 14'h2CBC;
            14'd 5861: out = 14'h2CBA;
            14'd 5862: out = 14'h2CB8;
            14'd 5863: out = 14'h2CB6;
            14'd 5864: out = 14'h2CB4;
            14'd 5865: out = 14'h2CB2;
            14'd 5866: out = 14'h2CB0;
            14'd 5867: out = 14'h2CAE;
            14'd 5868: out = 14'h2CAC;
            14'd 5869: out = 14'h2CAA;
            14'd 5870: out = 14'h2CA9;
            14'd 5871: out = 14'h2CA7;
            14'd 5872: out = 14'h2CA5;
            14'd 5873: out = 14'h2CA3;
            14'd 5874: out = 14'h2CA1;
            14'd 5875: out = 14'h2C9F;
            14'd 5876: out = 14'h2C9D;
            14'd 5877: out = 14'h2C9B;
            14'd 5878: out = 14'h2C99;
            14'd 5879: out = 14'h2C97;
            14'd 5880: out = 14'h2C95;
            14'd 5881: out = 14'h2C93;
            14'd 5882: out = 14'h2C91;
            14'd 5883: out = 14'h2C8F;
            14'd 5884: out = 14'h2C8D;
            14'd 5885: out = 14'h2C8B;
            14'd 5886: out = 14'h2C89;
            14'd 5887: out = 14'h2C88;
            14'd 5888: out = 14'h2C86;
            14'd 5889: out = 14'h2C84;
            14'd 5890: out = 14'h2C82;
            14'd 5891: out = 14'h2C80;
            14'd 5892: out = 14'h2C7E;
            14'd 5893: out = 14'h2C7C;
            14'd 5894: out = 14'h2C7A;
            14'd 5895: out = 14'h2C78;
            14'd 5896: out = 14'h2C76;
            14'd 5897: out = 14'h2C74;
            14'd 5898: out = 14'h2C72;
            14'd 5899: out = 14'h2C70;
            14'd 5900: out = 14'h2C6E;
            14'd 5901: out = 14'h2C6C;
            14'd 5902: out = 14'h2C6B;
            14'd 5903: out = 14'h2C69;
            14'd 5904: out = 14'h2C67;
            14'd 5905: out = 14'h2C65;
            14'd 5906: out = 14'h2C63;
            14'd 5907: out = 14'h2C61;
            14'd 5908: out = 14'h2C5F;
            14'd 5909: out = 14'h2C5D;
            14'd 5910: out = 14'h2C5B;
            14'd 5911: out = 14'h2C59;
            14'd 5912: out = 14'h2C57;
            14'd 5913: out = 14'h2C55;
            14'd 5914: out = 14'h2C53;
            14'd 5915: out = 14'h2C52;
            14'd 5916: out = 14'h2C50;
            14'd 5917: out = 14'h2C4E;
            14'd 5918: out = 14'h2C4C;
            14'd 5919: out = 14'h2C4A;
            14'd 5920: out = 14'h2C48;
            14'd 5921: out = 14'h2C46;
            14'd 5922: out = 14'h2C44;
            14'd 5923: out = 14'h2C42;
            14'd 5924: out = 14'h2C40;
            14'd 5925: out = 14'h2C3E;
            14'd 5926: out = 14'h2C3C;
            14'd 5927: out = 14'h2C3B;
            14'd 5928: out = 14'h2C39;
            14'd 5929: out = 14'h2C37;
            14'd 5930: out = 14'h2C35;
            14'd 5931: out = 14'h2C33;
            14'd 5932: out = 14'h2C31;
            14'd 5933: out = 14'h2C2F;
            14'd 5934: out = 14'h2C2D;
            14'd 5935: out = 14'h2C2B;
            14'd 5936: out = 14'h2C29;
            14'd 5937: out = 14'h2C27;
            14'd 5938: out = 14'h2C26;
            14'd 5939: out = 14'h2C24;
            14'd 5940: out = 14'h2C22;
            14'd 5941: out = 14'h2C20;
            14'd 5942: out = 14'h2C1E;
            14'd 5943: out = 14'h2C1C;
            14'd 5944: out = 14'h2C1A;
            14'd 5945: out = 14'h2C18;
            14'd 5946: out = 14'h2C16;
            14'd 5947: out = 14'h2C14;
            14'd 5948: out = 14'h2C13;
            14'd 5949: out = 14'h2C11;
            14'd 5950: out = 14'h2C0F;
            14'd 5951: out = 14'h2C0D;
            14'd 5952: out = 14'h2C0B;
            14'd 5953: out = 14'h2C09;
            14'd 5954: out = 14'h2C07;
            14'd 5955: out = 14'h2C05;
            14'd 5956: out = 14'h2C03;
            14'd 5957: out = 14'h2C02;
            14'd 5958: out = 14'h2C00;
            14'd 5959: out = 14'h2BFE;
            14'd 5960: out = 14'h2BFC;
            14'd 5961: out = 14'h2BFA;
            14'd 5962: out = 14'h2BF8;
            14'd 5963: out = 14'h2BF6;
            14'd 5964: out = 14'h2BF4;
            14'd 5965: out = 14'h2BF2;
            14'd 5966: out = 14'h2BF1;
            14'd 5967: out = 14'h2BEF;
            14'd 5968: out = 14'h2BED;
            14'd 5969: out = 14'h2BEB;
            14'd 5970: out = 14'h2BE9;
            14'd 5971: out = 14'h2BE7;
            14'd 5972: out = 14'h2BE5;
            14'd 5973: out = 14'h2BE3;
            14'd 5974: out = 14'h2BE1;
            14'd 5975: out = 14'h2BE0;
            14'd 5976: out = 14'h2BDE;
            14'd 5977: out = 14'h2BDC;
            14'd 5978: out = 14'h2BDA;
            14'd 5979: out = 14'h2BD8;
            14'd 5980: out = 14'h2BD6;
            14'd 5981: out = 14'h2BD4;
            14'd 5982: out = 14'h2BD2;
            14'd 5983: out = 14'h2BD1;
            14'd 5984: out = 14'h2BCF;
            14'd 5985: out = 14'h2BCD;
            14'd 5986: out = 14'h2BCB;
            14'd 5987: out = 14'h2BC9;
            14'd 5988: out = 14'h2BC7;
            14'd 5989: out = 14'h2BC5;
            14'd 5990: out = 14'h2BC3;
            14'd 5991: out = 14'h2BC2;
            14'd 5992: out = 14'h2BC0;
            14'd 5993: out = 14'h2BBE;
            14'd 5994: out = 14'h2BBC;
            14'd 5995: out = 14'h2BBA;
            14'd 5996: out = 14'h2BB8;
            14'd 5997: out = 14'h2BB6;
            14'd 5998: out = 14'h2BB5;
            14'd 5999: out = 14'h2BB3;
            14'd 6000: out = 14'h2BB1;
            14'd 6001: out = 14'h2BAF;
            14'd 6002: out = 14'h2BAD;
            14'd 6003: out = 14'h2BAB;
            14'd 6004: out = 14'h2BA9;
            14'd 6005: out = 14'h2BA7;
            14'd 6006: out = 14'h2BA6;
            14'd 6007: out = 14'h2BA4;
            14'd 6008: out = 14'h2BA2;
            14'd 6009: out = 14'h2BA0;
            14'd 6010: out = 14'h2B9E;
            14'd 6011: out = 14'h2B9C;
            14'd 6012: out = 14'h2B9A;
            14'd 6013: out = 14'h2B99;
            14'd 6014: out = 14'h2B97;
            14'd 6015: out = 14'h2B95;
            14'd 6016: out = 14'h2B93;
            14'd 6017: out = 14'h2B91;
            14'd 6018: out = 14'h2B8F;
            14'd 6019: out = 14'h2B8E;
            14'd 6020: out = 14'h2B8C;
            14'd 6021: out = 14'h2B8A;
            14'd 6022: out = 14'h2B88;
            14'd 6023: out = 14'h2B86;
            14'd 6024: out = 14'h2B84;
            14'd 6025: out = 14'h2B82;
            14'd 6026: out = 14'h2B81;
            14'd 6027: out = 14'h2B7F;
            14'd 6028: out = 14'h2B7D;
            14'd 6029: out = 14'h2B7B;
            14'd 6030: out = 14'h2B79;
            14'd 6031: out = 14'h2B77;
            14'd 6032: out = 14'h2B75;
            14'd 6033: out = 14'h2B74;
            14'd 6034: out = 14'h2B72;
            14'd 6035: out = 14'h2B70;
            14'd 6036: out = 14'h2B6E;
            14'd 6037: out = 14'h2B6C;
            14'd 6038: out = 14'h2B6A;
            14'd 6039: out = 14'h2B69;
            14'd 6040: out = 14'h2B67;
            14'd 6041: out = 14'h2B65;
            14'd 6042: out = 14'h2B63;
            14'd 6043: out = 14'h2B61;
            14'd 6044: out = 14'h2B5F;
            14'd 6045: out = 14'h2B5E;
            14'd 6046: out = 14'h2B5C;
            14'd 6047: out = 14'h2B5A;
            14'd 6048: out = 14'h2B58;
            14'd 6049: out = 14'h2B56;
            14'd 6050: out = 14'h2B54;
            14'd 6051: out = 14'h2B53;
            14'd 6052: out = 14'h2B51;
            14'd 6053: out = 14'h2B4F;
            14'd 6054: out = 14'h2B4D;
            14'd 6055: out = 14'h2B4B;
            14'd 6056: out = 14'h2B49;
            14'd 6057: out = 14'h2B48;
            14'd 6058: out = 14'h2B46;
            14'd 6059: out = 14'h2B44;
            14'd 6060: out = 14'h2B42;
            14'd 6061: out = 14'h2B40;
            14'd 6062: out = 14'h2B3E;
            14'd 6063: out = 14'h2B3D;
            14'd 6064: out = 14'h2B3B;
            14'd 6065: out = 14'h2B39;
            14'd 6066: out = 14'h2B37;
            14'd 6067: out = 14'h2B35;
            14'd 6068: out = 14'h2B33;
            14'd 6069: out = 14'h2B32;
            14'd 6070: out = 14'h2B30;
            14'd 6071: out = 14'h2B2E;
            14'd 6072: out = 14'h2B2C;
            14'd 6073: out = 14'h2B2A;
            14'd 6074: out = 14'h2B29;
            14'd 6075: out = 14'h2B27;
            14'd 6076: out = 14'h2B25;
            14'd 6077: out = 14'h2B23;
            14'd 6078: out = 14'h2B21;
            14'd 6079: out = 14'h2B1F;
            14'd 6080: out = 14'h2B1E;
            14'd 6081: out = 14'h2B1C;
            14'd 6082: out = 14'h2B1A;
            14'd 6083: out = 14'h2B18;
            14'd 6084: out = 14'h2B16;
            14'd 6085: out = 14'h2B15;
            14'd 6086: out = 14'h2B13;
            14'd 6087: out = 14'h2B11;
            14'd 6088: out = 14'h2B0F;
            14'd 6089: out = 14'h2B0D;
            14'd 6090: out = 14'h2B0C;
            14'd 6091: out = 14'h2B0A;
            14'd 6092: out = 14'h2B08;
            14'd 6093: out = 14'h2B06;
            14'd 6094: out = 14'h2B04;
            14'd 6095: out = 14'h2B02;
            14'd 6096: out = 14'h2B01;
            14'd 6097: out = 14'h2AFF;
            14'd 6098: out = 14'h2AFD;
            14'd 6099: out = 14'h2AFB;
            14'd 6100: out = 14'h2AF9;
            14'd 6101: out = 14'h2AF8;
            14'd 6102: out = 14'h2AF6;
            14'd 6103: out = 14'h2AF4;
            14'd 6104: out = 14'h2AF2;
            14'd 6105: out = 14'h2AF0;
            14'd 6106: out = 14'h2AEF;
            14'd 6107: out = 14'h2AED;
            14'd 6108: out = 14'h2AEB;
            14'd 6109: out = 14'h2AE9;
            14'd 6110: out = 14'h2AE7;
            14'd 6111: out = 14'h2AE6;
            14'd 6112: out = 14'h2AE4;
            14'd 6113: out = 14'h2AE2;
            14'd 6114: out = 14'h2AE0;
            14'd 6115: out = 14'h2ADE;
            14'd 6116: out = 14'h2ADD;
            14'd 6117: out = 14'h2ADB;
            14'd 6118: out = 14'h2AD9;
            14'd 6119: out = 14'h2AD7;
            14'd 6120: out = 14'h2AD6;
            14'd 6121: out = 14'h2AD4;
            14'd 6122: out = 14'h2AD2;
            14'd 6123: out = 14'h2AD0;
            14'd 6124: out = 14'h2ACE;
            14'd 6125: out = 14'h2ACD;
            14'd 6126: out = 14'h2ACB;
            14'd 6127: out = 14'h2AC9;
            14'd 6128: out = 14'h2AC7;
            14'd 6129: out = 14'h2AC5;
            14'd 6130: out = 14'h2AC4;
            14'd 6131: out = 14'h2AC2;
            14'd 6132: out = 14'h2AC0;
            14'd 6133: out = 14'h2ABE;
            14'd 6134: out = 14'h2ABC;
            14'd 6135: out = 14'h2ABB;
            14'd 6136: out = 14'h2AB9;
            14'd 6137: out = 14'h2AB7;
            14'd 6138: out = 14'h2AB5;
            14'd 6139: out = 14'h2AB4;
            14'd 6140: out = 14'h2AB2;
            14'd 6141: out = 14'h2AB0;
            14'd 6142: out = 14'h2AAE;
            14'd 6143: out = 14'h2AAC;
            14'd 6144: out = 14'h2AAB;
            14'd 6145: out = 14'h2AA9;
            14'd 6146: out = 14'h2AA7;
            14'd 6147: out = 14'h2AA5;
            14'd 6148: out = 14'h2AA4;
            14'd 6149: out = 14'h2AA2;
            14'd 6150: out = 14'h2AA0;
            14'd 6151: out = 14'h2A9E;
            14'd 6152: out = 14'h2A9C;
            14'd 6153: out = 14'h2A9B;
            14'd 6154: out = 14'h2A99;
            14'd 6155: out = 14'h2A97;
            14'd 6156: out = 14'h2A95;
            14'd 6157: out = 14'h2A94;
            14'd 6158: out = 14'h2A92;
            14'd 6159: out = 14'h2A90;
            14'd 6160: out = 14'h2A8E;
            14'd 6161: out = 14'h2A8D;
            14'd 6162: out = 14'h2A8B;
            14'd 6163: out = 14'h2A89;
            14'd 6164: out = 14'h2A87;
            14'd 6165: out = 14'h2A85;
            14'd 6166: out = 14'h2A84;
            14'd 6167: out = 14'h2A82;
            14'd 6168: out = 14'h2A80;
            14'd 6169: out = 14'h2A7E;
            14'd 6170: out = 14'h2A7D;
            14'd 6171: out = 14'h2A7B;
            14'd 6172: out = 14'h2A79;
            14'd 6173: out = 14'h2A77;
            14'd 6174: out = 14'h2A76;
            14'd 6175: out = 14'h2A74;
            14'd 6176: out = 14'h2A72;
            14'd 6177: out = 14'h2A70;
            14'd 6178: out = 14'h2A6F;
            14'd 6179: out = 14'h2A6D;
            14'd 6180: out = 14'h2A6B;
            14'd 6181: out = 14'h2A69;
            14'd 6182: out = 14'h2A68;
            14'd 6183: out = 14'h2A66;
            14'd 6184: out = 14'h2A64;
            14'd 6185: out = 14'h2A62;
            14'd 6186: out = 14'h2A61;
            14'd 6187: out = 14'h2A5F;
            14'd 6188: out = 14'h2A5D;
            14'd 6189: out = 14'h2A5B;
            14'd 6190: out = 14'h2A59;
            14'd 6191: out = 14'h2A58;
            14'd 6192: out = 14'h2A56;
            14'd 6193: out = 14'h2A54;
            14'd 6194: out = 14'h2A52;
            14'd 6195: out = 14'h2A51;
            14'd 6196: out = 14'h2A4F;
            14'd 6197: out = 14'h2A4D;
            14'd 6198: out = 14'h2A4C;
            14'd 6199: out = 14'h2A4A;
            14'd 6200: out = 14'h2A48;
            14'd 6201: out = 14'h2A46;
            14'd 6202: out = 14'h2A45;
            14'd 6203: out = 14'h2A43;
            14'd 6204: out = 14'h2A41;
            14'd 6205: out = 14'h2A3F;
            14'd 6206: out = 14'h2A3E;
            14'd 6207: out = 14'h2A3C;
            14'd 6208: out = 14'h2A3A;
            14'd 6209: out = 14'h2A38;
            14'd 6210: out = 14'h2A37;
            14'd 6211: out = 14'h2A35;
            14'd 6212: out = 14'h2A33;
            14'd 6213: out = 14'h2A31;
            14'd 6214: out = 14'h2A30;
            14'd 6215: out = 14'h2A2E;
            14'd 6216: out = 14'h2A2C;
            14'd 6217: out = 14'h2A2A;
            14'd 6218: out = 14'h2A29;
            14'd 6219: out = 14'h2A27;
            14'd 6220: out = 14'h2A25;
            14'd 6221: out = 14'h2A23;
            14'd 6222: out = 14'h2A22;
            14'd 6223: out = 14'h2A20;
            14'd 6224: out = 14'h2A1E;
            14'd 6225: out = 14'h2A1D;
            14'd 6226: out = 14'h2A1B;
            14'd 6227: out = 14'h2A19;
            14'd 6228: out = 14'h2A17;
            14'd 6229: out = 14'h2A16;
            14'd 6230: out = 14'h2A14;
            14'd 6231: out = 14'h2A12;
            14'd 6232: out = 14'h2A10;
            14'd 6233: out = 14'h2A0F;
            14'd 6234: out = 14'h2A0D;
            14'd 6235: out = 14'h2A0B;
            14'd 6236: out = 14'h2A0A;
            14'd 6237: out = 14'h2A08;
            14'd 6238: out = 14'h2A06;
            14'd 6239: out = 14'h2A04;
            14'd 6240: out = 14'h2A03;
            14'd 6241: out = 14'h2A01;
            14'd 6242: out = 14'h29FF;
            14'd 6243: out = 14'h29FD;
            14'd 6244: out = 14'h29FC;
            14'd 6245: out = 14'h29FA;
            14'd 6246: out = 14'h29F8;
            14'd 6247: out = 14'h29F7;
            14'd 6248: out = 14'h29F5;
            14'd 6249: out = 14'h29F3;
            14'd 6250: out = 14'h29F1;
            14'd 6251: out = 14'h29F0;
            14'd 6252: out = 14'h29EE;
            14'd 6253: out = 14'h29EC;
            14'd 6254: out = 14'h29EB;
            14'd 6255: out = 14'h29E9;
            14'd 6256: out = 14'h29E7;
            14'd 6257: out = 14'h29E5;
            14'd 6258: out = 14'h29E4;
            14'd 6259: out = 14'h29E2;
            14'd 6260: out = 14'h29E0;
            14'd 6261: out = 14'h29DF;
            14'd 6262: out = 14'h29DD;
            14'd 6263: out = 14'h29DB;
            14'd 6264: out = 14'h29D9;
            14'd 6265: out = 14'h29D8;
            14'd 6266: out = 14'h29D6;
            14'd 6267: out = 14'h29D4;
            14'd 6268: out = 14'h29D3;
            14'd 6269: out = 14'h29D1;
            14'd 6270: out = 14'h29CF;
            14'd 6271: out = 14'h29CD;
            14'd 6272: out = 14'h29CC;
            14'd 6273: out = 14'h29CA;
            14'd 6274: out = 14'h29C8;
            14'd 6275: out = 14'h29C7;
            14'd 6276: out = 14'h29C5;
            14'd 6277: out = 14'h29C3;
            14'd 6278: out = 14'h29C2;
            14'd 6279: out = 14'h29C0;
            14'd 6280: out = 14'h29BE;
            14'd 6281: out = 14'h29BC;
            14'd 6282: out = 14'h29BB;
            14'd 6283: out = 14'h29B9;
            14'd 6284: out = 14'h29B7;
            14'd 6285: out = 14'h29B6;
            14'd 6286: out = 14'h29B4;
            14'd 6287: out = 14'h29B2;
            14'd 6288: out = 14'h29B1;
            14'd 6289: out = 14'h29AF;
            14'd 6290: out = 14'h29AD;
            14'd 6291: out = 14'h29AB;
            14'd 6292: out = 14'h29AA;
            14'd 6293: out = 14'h29A8;
            14'd 6294: out = 14'h29A6;
            14'd 6295: out = 14'h29A5;
            14'd 6296: out = 14'h29A3;
            14'd 6297: out = 14'h29A1;
            14'd 6298: out = 14'h29A0;
            14'd 6299: out = 14'h299E;
            14'd 6300: out = 14'h299C;
            14'd 6301: out = 14'h299B;
            14'd 6302: out = 14'h2999;
            14'd 6303: out = 14'h2997;
            14'd 6304: out = 14'h2995;
            14'd 6305: out = 14'h2994;
            14'd 6306: out = 14'h2992;
            14'd 6307: out = 14'h2990;
            14'd 6308: out = 14'h298F;
            14'd 6309: out = 14'h298D;
            14'd 6310: out = 14'h298B;
            14'd 6311: out = 14'h298A;
            14'd 6312: out = 14'h2988;
            14'd 6313: out = 14'h2986;
            14'd 6314: out = 14'h2985;
            14'd 6315: out = 14'h2983;
            14'd 6316: out = 14'h2981;
            14'd 6317: out = 14'h2980;
            14'd 6318: out = 14'h297E;
            14'd 6319: out = 14'h297C;
            14'd 6320: out = 14'h297A;
            14'd 6321: out = 14'h2979;
            14'd 6322: out = 14'h2977;
            14'd 6323: out = 14'h2975;
            14'd 6324: out = 14'h2974;
            14'd 6325: out = 14'h2972;
            14'd 6326: out = 14'h2970;
            14'd 6327: out = 14'h296F;
            14'd 6328: out = 14'h296D;
            14'd 6329: out = 14'h296B;
            14'd 6330: out = 14'h296A;
            14'd 6331: out = 14'h2968;
            14'd 6332: out = 14'h2966;
            14'd 6333: out = 14'h2965;
            14'd 6334: out = 14'h2963;
            14'd 6335: out = 14'h2961;
            14'd 6336: out = 14'h2960;
            14'd 6337: out = 14'h295E;
            14'd 6338: out = 14'h295C;
            14'd 6339: out = 14'h295B;
            14'd 6340: out = 14'h2959;
            14'd 6341: out = 14'h2957;
            14'd 6342: out = 14'h2956;
            14'd 6343: out = 14'h2954;
            14'd 6344: out = 14'h2952;
            14'd 6345: out = 14'h2951;
            14'd 6346: out = 14'h294F;
            14'd 6347: out = 14'h294D;
            14'd 6348: out = 14'h294C;
            14'd 6349: out = 14'h294A;
            14'd 6350: out = 14'h2948;
            14'd 6351: out = 14'h2947;
            14'd 6352: out = 14'h2945;
            14'd 6353: out = 14'h2943;
            14'd 6354: out = 14'h2942;
            14'd 6355: out = 14'h2940;
            14'd 6356: out = 14'h293E;
            14'd 6357: out = 14'h293D;
            14'd 6358: out = 14'h293B;
            14'd 6359: out = 14'h2939;
            14'd 6360: out = 14'h2938;
            14'd 6361: out = 14'h2936;
            14'd 6362: out = 14'h2934;
            14'd 6363: out = 14'h2933;
            14'd 6364: out = 14'h2931;
            14'd 6365: out = 14'h292F;
            14'd 6366: out = 14'h292E;
            14'd 6367: out = 14'h292C;
            14'd 6368: out = 14'h292A;
            14'd 6369: out = 14'h2929;
            14'd 6370: out = 14'h2927;
            14'd 6371: out = 14'h2925;
            14'd 6372: out = 14'h2924;
            14'd 6373: out = 14'h2922;
            14'd 6374: out = 14'h2921;
            14'd 6375: out = 14'h291F;
            14'd 6376: out = 14'h291D;
            14'd 6377: out = 14'h291C;
            14'd 6378: out = 14'h291A;
            14'd 6379: out = 14'h2918;
            14'd 6380: out = 14'h2917;
            14'd 6381: out = 14'h2915;
            14'd 6382: out = 14'h2913;
            14'd 6383: out = 14'h2912;
            14'd 6384: out = 14'h2910;
            14'd 6385: out = 14'h290E;
            14'd 6386: out = 14'h290D;
            14'd 6387: out = 14'h290B;
            14'd 6388: out = 14'h2909;
            14'd 6389: out = 14'h2908;
            14'd 6390: out = 14'h2906;
            14'd 6391: out = 14'h2905;
            14'd 6392: out = 14'h2903;
            14'd 6393: out = 14'h2901;
            14'd 6394: out = 14'h2900;
            14'd 6395: out = 14'h28FE;
            14'd 6396: out = 14'h28FC;
            14'd 6397: out = 14'h28FB;
            14'd 6398: out = 14'h28F9;
            14'd 6399: out = 14'h28F7;
            14'd 6400: out = 14'h28F6;
            14'd 6401: out = 14'h28F4;
            14'd 6402: out = 14'h28F2;
            14'd 6403: out = 14'h28F1;
            14'd 6404: out = 14'h28EF;
            14'd 6405: out = 14'h28EE;
            14'd 6406: out = 14'h28EC;
            14'd 6407: out = 14'h28EA;
            14'd 6408: out = 14'h28E9;
            14'd 6409: out = 14'h28E7;
            14'd 6410: out = 14'h28E5;
            14'd 6411: out = 14'h28E4;
            14'd 6412: out = 14'h28E2;
            14'd 6413: out = 14'h28E1;
            14'd 6414: out = 14'h28DF;
            14'd 6415: out = 14'h28DD;
            14'd 6416: out = 14'h28DC;
            14'd 6417: out = 14'h28DA;
            14'd 6418: out = 14'h28D8;
            14'd 6419: out = 14'h28D7;
            14'd 6420: out = 14'h28D5;
            14'd 6421: out = 14'h28D3;
            14'd 6422: out = 14'h28D2;
            14'd 6423: out = 14'h28D0;
            14'd 6424: out = 14'h28CF;
            14'd 6425: out = 14'h28CD;
            14'd 6426: out = 14'h28CB;
            14'd 6427: out = 14'h28CA;
            14'd 6428: out = 14'h28C8;
            14'd 6429: out = 14'h28C6;
            14'd 6430: out = 14'h28C5;
            14'd 6431: out = 14'h28C3;
            14'd 6432: out = 14'h28C2;
            14'd 6433: out = 14'h28C0;
            14'd 6434: out = 14'h28BE;
            14'd 6435: out = 14'h28BD;
            14'd 6436: out = 14'h28BB;
            14'd 6437: out = 14'h28B9;
            14'd 6438: out = 14'h28B8;
            14'd 6439: out = 14'h28B6;
            14'd 6440: out = 14'h28B5;
            14'd 6441: out = 14'h28B3;
            14'd 6442: out = 14'h28B1;
            14'd 6443: out = 14'h28B0;
            14'd 6444: out = 14'h28AE;
            14'd 6445: out = 14'h28AD;
            14'd 6446: out = 14'h28AB;
            14'd 6447: out = 14'h28A9;
            14'd 6448: out = 14'h28A8;
            14'd 6449: out = 14'h28A6;
            14'd 6450: out = 14'h28A4;
            14'd 6451: out = 14'h28A3;
            14'd 6452: out = 14'h28A1;
            14'd 6453: out = 14'h28A0;
            14'd 6454: out = 14'h289E;
            14'd 6455: out = 14'h289C;
            14'd 6456: out = 14'h289B;
            14'd 6457: out = 14'h2899;
            14'd 6458: out = 14'h2898;
            14'd 6459: out = 14'h2896;
            14'd 6460: out = 14'h2894;
            14'd 6461: out = 14'h2893;
            14'd 6462: out = 14'h2891;
            14'd 6463: out = 14'h2890;
            14'd 6464: out = 14'h288E;
            14'd 6465: out = 14'h288C;
            14'd 6466: out = 14'h288B;
            14'd 6467: out = 14'h2889;
            14'd 6468: out = 14'h2888;
            14'd 6469: out = 14'h2886;
            14'd 6470: out = 14'h2884;
            14'd 6471: out = 14'h2883;
            14'd 6472: out = 14'h2881;
            14'd 6473: out = 14'h2880;
            14'd 6474: out = 14'h287E;
            14'd 6475: out = 14'h287C;
            14'd 6476: out = 14'h287B;
            14'd 6477: out = 14'h2879;
            14'd 6478: out = 14'h2878;
            14'd 6479: out = 14'h2876;
            14'd 6480: out = 14'h2874;
            14'd 6481: out = 14'h2873;
            14'd 6482: out = 14'h2871;
            14'd 6483: out = 14'h2870;
            14'd 6484: out = 14'h286E;
            14'd 6485: out = 14'h286C;
            14'd 6486: out = 14'h286B;
            14'd 6487: out = 14'h2869;
            14'd 6488: out = 14'h2868;
            14'd 6489: out = 14'h2866;
            14'd 6490: out = 14'h2864;
            14'd 6491: out = 14'h2863;
            14'd 6492: out = 14'h2861;
            14'd 6493: out = 14'h2860;
            14'd 6494: out = 14'h285E;
            14'd 6495: out = 14'h285C;
            14'd 6496: out = 14'h285B;
            14'd 6497: out = 14'h2859;
            14'd 6498: out = 14'h2858;
            14'd 6499: out = 14'h2856;
            14'd 6500: out = 14'h2854;
            14'd 6501: out = 14'h2853;
            14'd 6502: out = 14'h2851;
            14'd 6503: out = 14'h2850;
            14'd 6504: out = 14'h284E;
            14'd 6505: out = 14'h284D;
            14'd 6506: out = 14'h284B;
            14'd 6507: out = 14'h2849;
            14'd 6508: out = 14'h2848;
            14'd 6509: out = 14'h2846;
            14'd 6510: out = 14'h2845;
            14'd 6511: out = 14'h2843;
            14'd 6512: out = 14'h2841;
            14'd 6513: out = 14'h2840;
            14'd 6514: out = 14'h283E;
            14'd 6515: out = 14'h283D;
            14'd 6516: out = 14'h283B;
            14'd 6517: out = 14'h283A;
            14'd 6518: out = 14'h2838;
            14'd 6519: out = 14'h2836;
            14'd 6520: out = 14'h2835;
            14'd 6521: out = 14'h2833;
            14'd 6522: out = 14'h2832;
            14'd 6523: out = 14'h2830;
            14'd 6524: out = 14'h282E;
            14'd 6525: out = 14'h282D;
            14'd 6526: out = 14'h282B;
            14'd 6527: out = 14'h282A;
            14'd 6528: out = 14'h2828;
            14'd 6529: out = 14'h2827;
            14'd 6530: out = 14'h2825;
            14'd 6531: out = 14'h2823;
            14'd 6532: out = 14'h2822;
            14'd 6533: out = 14'h2820;
            14'd 6534: out = 14'h281F;
            14'd 6535: out = 14'h281D;
            14'd 6536: out = 14'h281C;
            14'd 6537: out = 14'h281A;
            14'd 6538: out = 14'h2818;
            14'd 6539: out = 14'h2817;
            14'd 6540: out = 14'h2815;
            14'd 6541: out = 14'h2814;
            14'd 6542: out = 14'h2812;
            14'd 6543: out = 14'h2811;
            14'd 6544: out = 14'h280F;
            14'd 6545: out = 14'h280D;
            14'd 6546: out = 14'h280C;
            14'd 6547: out = 14'h280A;
            14'd 6548: out = 14'h2809;
            14'd 6549: out = 14'h2807;
            14'd 6550: out = 14'h2806;
            14'd 6551: out = 14'h2804;
            14'd 6552: out = 14'h2803;
            14'd 6553: out = 14'h2801;
            14'd 6554: out = 14'h27FF;
            14'd 6555: out = 14'h27FE;
            14'd 6556: out = 14'h27FC;
            14'd 6557: out = 14'h27FB;
            14'd 6558: out = 14'h27F9;
            14'd 6559: out = 14'h27F8;
            14'd 6560: out = 14'h27F6;
            14'd 6561: out = 14'h27F4;
            14'd 6562: out = 14'h27F3;
            14'd 6563: out = 14'h27F1;
            14'd 6564: out = 14'h27F0;
            14'd 6565: out = 14'h27EE;
            14'd 6566: out = 14'h27ED;
            14'd 6567: out = 14'h27EB;
            14'd 6568: out = 14'h27EA;
            14'd 6569: out = 14'h27E8;
            14'd 6570: out = 14'h27E6;
            14'd 6571: out = 14'h27E5;
            14'd 6572: out = 14'h27E3;
            14'd 6573: out = 14'h27E2;
            14'd 6574: out = 14'h27E0;
            14'd 6575: out = 14'h27DF;
            14'd 6576: out = 14'h27DD;
            14'd 6577: out = 14'h27DC;
            14'd 6578: out = 14'h27DA;
            14'd 6579: out = 14'h27D8;
            14'd 6580: out = 14'h27D7;
            14'd 6581: out = 14'h27D5;
            14'd 6582: out = 14'h27D4;
            14'd 6583: out = 14'h27D2;
            14'd 6584: out = 14'h27D1;
            14'd 6585: out = 14'h27CF;
            14'd 6586: out = 14'h27CE;
            14'd 6587: out = 14'h27CC;
            14'd 6588: out = 14'h27CB;
            14'd 6589: out = 14'h27C9;
            14'd 6590: out = 14'h27C7;
            14'd 6591: out = 14'h27C6;
            14'd 6592: out = 14'h27C4;
            14'd 6593: out = 14'h27C3;
            14'd 6594: out = 14'h27C1;
            14'd 6595: out = 14'h27C0;
            14'd 6596: out = 14'h27BE;
            14'd 6597: out = 14'h27BD;
            14'd 6598: out = 14'h27BB;
            14'd 6599: out = 14'h27BA;
            14'd 6600: out = 14'h27B8;
            14'd 6601: out = 14'h27B6;
            14'd 6602: out = 14'h27B5;
            14'd 6603: out = 14'h27B3;
            14'd 6604: out = 14'h27B2;
            14'd 6605: out = 14'h27B0;
            14'd 6606: out = 14'h27AF;
            14'd 6607: out = 14'h27AD;
            14'd 6608: out = 14'h27AC;
            14'd 6609: out = 14'h27AA;
            14'd 6610: out = 14'h27A9;
            14'd 6611: out = 14'h27A7;
            14'd 6612: out = 14'h27A6;
            14'd 6613: out = 14'h27A4;
            14'd 6614: out = 14'h27A2;
            14'd 6615: out = 14'h27A1;
            14'd 6616: out = 14'h279F;
            14'd 6617: out = 14'h279E;
            14'd 6618: out = 14'h279C;
            14'd 6619: out = 14'h279B;
            14'd 6620: out = 14'h2799;
            14'd 6621: out = 14'h2798;
            14'd 6622: out = 14'h2796;
            14'd 6623: out = 14'h2795;
            14'd 6624: out = 14'h2793;
            14'd 6625: out = 14'h2792;
            14'd 6626: out = 14'h2790;
            14'd 6627: out = 14'h278F;
            14'd 6628: out = 14'h278D;
            14'd 6629: out = 14'h278C;
            14'd 6630: out = 14'h278A;
            14'd 6631: out = 14'h2788;
            14'd 6632: out = 14'h2787;
            14'd 6633: out = 14'h2785;
            14'd 6634: out = 14'h2784;
            14'd 6635: out = 14'h2782;
            14'd 6636: out = 14'h2781;
            14'd 6637: out = 14'h277F;
            14'd 6638: out = 14'h277E;
            14'd 6639: out = 14'h277C;
            14'd 6640: out = 14'h277B;
            14'd 6641: out = 14'h2779;
            14'd 6642: out = 14'h2778;
            14'd 6643: out = 14'h2776;
            14'd 6644: out = 14'h2775;
            14'd 6645: out = 14'h2773;
            14'd 6646: out = 14'h2772;
            14'd 6647: out = 14'h2770;
            14'd 6648: out = 14'h276F;
            14'd 6649: out = 14'h276D;
            14'd 6650: out = 14'h276C;
            14'd 6651: out = 14'h276A;
            14'd 6652: out = 14'h2769;
            14'd 6653: out = 14'h2767;
            14'd 6654: out = 14'h2765;
            14'd 6655: out = 14'h2764;
            14'd 6656: out = 14'h2762;
            14'd 6657: out = 14'h2761;
            14'd 6658: out = 14'h275F;
            14'd 6659: out = 14'h275E;
            14'd 6660: out = 14'h275C;
            14'd 6661: out = 14'h275B;
            14'd 6662: out = 14'h2759;
            14'd 6663: out = 14'h2758;
            14'd 6664: out = 14'h2756;
            14'd 6665: out = 14'h2755;
            14'd 6666: out = 14'h2753;
            14'd 6667: out = 14'h2752;
            14'd 6668: out = 14'h2750;
            14'd 6669: out = 14'h274F;
            14'd 6670: out = 14'h274D;
            14'd 6671: out = 14'h274C;
            14'd 6672: out = 14'h274A;
            14'd 6673: out = 14'h2749;
            14'd 6674: out = 14'h2747;
            14'd 6675: out = 14'h2746;
            14'd 6676: out = 14'h2744;
            14'd 6677: out = 14'h2743;
            14'd 6678: out = 14'h2741;
            14'd 6679: out = 14'h2740;
            14'd 6680: out = 14'h273E;
            14'd 6681: out = 14'h273D;
            14'd 6682: out = 14'h273B;
            14'd 6683: out = 14'h273A;
            14'd 6684: out = 14'h2738;
            14'd 6685: out = 14'h2737;
            14'd 6686: out = 14'h2735;
            14'd 6687: out = 14'h2734;
            14'd 6688: out = 14'h2732;
            14'd 6689: out = 14'h2731;
            14'd 6690: out = 14'h272F;
            14'd 6691: out = 14'h272E;
            14'd 6692: out = 14'h272C;
            14'd 6693: out = 14'h272B;
            14'd 6694: out = 14'h2729;
            14'd 6695: out = 14'h2728;
            14'd 6696: out = 14'h2726;
            14'd 6697: out = 14'h2725;
            14'd 6698: out = 14'h2723;
            14'd 6699: out = 14'h2722;
            14'd 6700: out = 14'h2720;
            14'd 6701: out = 14'h271F;
            14'd 6702: out = 14'h271D;
            14'd 6703: out = 14'h271C;
            14'd 6704: out = 14'h271A;
            14'd 6705: out = 14'h2719;
            14'd 6706: out = 14'h2717;
            14'd 6707: out = 14'h2716;
            14'd 6708: out = 14'h2714;
            14'd 6709: out = 14'h2713;
            14'd 6710: out = 14'h2711;
            14'd 6711: out = 14'h2710;
            14'd 6712: out = 14'h270E;
            14'd 6713: out = 14'h270D;
            14'd 6714: out = 14'h270B;
            14'd 6715: out = 14'h270A;
            14'd 6716: out = 14'h2708;
            14'd 6717: out = 14'h2707;
            14'd 6718: out = 14'h2705;
            14'd 6719: out = 14'h2704;
            14'd 6720: out = 14'h2702;
            14'd 6721: out = 14'h2701;
            14'd 6722: out = 14'h26FF;
            14'd 6723: out = 14'h26FE;
            14'd 6724: out = 14'h26FC;
            14'd 6725: out = 14'h26FB;
            14'd 6726: out = 14'h26FA;
            14'd 6727: out = 14'h26F8;
            14'd 6728: out = 14'h26F7;
            14'd 6729: out = 14'h26F5;
            14'd 6730: out = 14'h26F4;
            14'd 6731: out = 14'h26F2;
            14'd 6732: out = 14'h26F1;
            14'd 6733: out = 14'h26EF;
            14'd 6734: out = 14'h26EE;
            14'd 6735: out = 14'h26EC;
            14'd 6736: out = 14'h26EB;
            14'd 6737: out = 14'h26E9;
            14'd 6738: out = 14'h26E8;
            14'd 6739: out = 14'h26E6;
            14'd 6740: out = 14'h26E5;
            14'd 6741: out = 14'h26E3;
            14'd 6742: out = 14'h26E2;
            14'd 6743: out = 14'h26E0;
            14'd 6744: out = 14'h26DF;
            14'd 6745: out = 14'h26DD;
            14'd 6746: out = 14'h26DC;
            14'd 6747: out = 14'h26DA;
            14'd 6748: out = 14'h26D9;
            14'd 6749: out = 14'h26D8;
            14'd 6750: out = 14'h26D6;
            14'd 6751: out = 14'h26D5;
            14'd 6752: out = 14'h26D3;
            14'd 6753: out = 14'h26D2;
            14'd 6754: out = 14'h26D0;
            14'd 6755: out = 14'h26CF;
            14'd 6756: out = 14'h26CD;
            14'd 6757: out = 14'h26CC;
            14'd 6758: out = 14'h26CA;
            14'd 6759: out = 14'h26C9;
            14'd 6760: out = 14'h26C7;
            14'd 6761: out = 14'h26C6;
            14'd 6762: out = 14'h26C4;
            14'd 6763: out = 14'h26C3;
            14'd 6764: out = 14'h26C1;
            14'd 6765: out = 14'h26C0;
            14'd 6766: out = 14'h26BF;
            14'd 6767: out = 14'h26BD;
            14'd 6768: out = 14'h26BC;
            14'd 6769: out = 14'h26BA;
            14'd 6770: out = 14'h26B9;
            14'd 6771: out = 14'h26B7;
            14'd 6772: out = 14'h26B6;
            14'd 6773: out = 14'h26B4;
            14'd 6774: out = 14'h26B3;
            14'd 6775: out = 14'h26B1;
            14'd 6776: out = 14'h26B0;
            14'd 6777: out = 14'h26AE;
            14'd 6778: out = 14'h26AD;
            14'd 6779: out = 14'h26AC;
            14'd 6780: out = 14'h26AA;
            14'd 6781: out = 14'h26A9;
            14'd 6782: out = 14'h26A7;
            14'd 6783: out = 14'h26A6;
            14'd 6784: out = 14'h26A4;
            14'd 6785: out = 14'h26A3;
            14'd 6786: out = 14'h26A1;
            14'd 6787: out = 14'h26A0;
            14'd 6788: out = 14'h269E;
            14'd 6789: out = 14'h269D;
            14'd 6790: out = 14'h269B;
            14'd 6791: out = 14'h269A;
            14'd 6792: out = 14'h2699;
            14'd 6793: out = 14'h2697;
            14'd 6794: out = 14'h2696;
            14'd 6795: out = 14'h2694;
            14'd 6796: out = 14'h2693;
            14'd 6797: out = 14'h2691;
            14'd 6798: out = 14'h2690;
            14'd 6799: out = 14'h268E;
            14'd 6800: out = 14'h268D;
            14'd 6801: out = 14'h268B;
            14'd 6802: out = 14'h268A;
            14'd 6803: out = 14'h2689;
            14'd 6804: out = 14'h2687;
            14'd 6805: out = 14'h2686;
            14'd 6806: out = 14'h2684;
            14'd 6807: out = 14'h2683;
            14'd 6808: out = 14'h2681;
            14'd 6809: out = 14'h2680;
            14'd 6810: out = 14'h267E;
            14'd 6811: out = 14'h267D;
            14'd 6812: out = 14'h267C;
            14'd 6813: out = 14'h267A;
            14'd 6814: out = 14'h2679;
            14'd 6815: out = 14'h2677;
            14'd 6816: out = 14'h2676;
            14'd 6817: out = 14'h2674;
            14'd 6818: out = 14'h2673;
            14'd 6819: out = 14'h2671;
            14'd 6820: out = 14'h2670;
            14'd 6821: out = 14'h266F;
            14'd 6822: out = 14'h266D;
            14'd 6823: out = 14'h266C;
            14'd 6824: out = 14'h266A;
            14'd 6825: out = 14'h2669;
            14'd 6826: out = 14'h2667;
            14'd 6827: out = 14'h2666;
            14'd 6828: out = 14'h2664;
            14'd 6829: out = 14'h2663;
            14'd 6830: out = 14'h2662;
            14'd 6831: out = 14'h2660;
            14'd 6832: out = 14'h265F;
            14'd 6833: out = 14'h265D;
            14'd 6834: out = 14'h265C;
            14'd 6835: out = 14'h265A;
            14'd 6836: out = 14'h2659;
            14'd 6837: out = 14'h2658;
            14'd 6838: out = 14'h2656;
            14'd 6839: out = 14'h2655;
            14'd 6840: out = 14'h2653;
            14'd 6841: out = 14'h2652;
            14'd 6842: out = 14'h2650;
            14'd 6843: out = 14'h264F;
            14'd 6844: out = 14'h264E;
            14'd 6845: out = 14'h264C;
            14'd 6846: out = 14'h264B;
            14'd 6847: out = 14'h2649;
            14'd 6848: out = 14'h2648;
            14'd 6849: out = 14'h2646;
            14'd 6850: out = 14'h2645;
            14'd 6851: out = 14'h2643;
            14'd 6852: out = 14'h2642;
            14'd 6853: out = 14'h2641;
            14'd 6854: out = 14'h263F;
            14'd 6855: out = 14'h263E;
            14'd 6856: out = 14'h263C;
            14'd 6857: out = 14'h263B;
            14'd 6858: out = 14'h2639;
            14'd 6859: out = 14'h2638;
            14'd 6860: out = 14'h2637;
            14'd 6861: out = 14'h2635;
            14'd 6862: out = 14'h2634;
            14'd 6863: out = 14'h2632;
            14'd 6864: out = 14'h2631;
            14'd 6865: out = 14'h2630;
            14'd 6866: out = 14'h262E;
            14'd 6867: out = 14'h262D;
            14'd 6868: out = 14'h262B;
            14'd 6869: out = 14'h262A;
            14'd 6870: out = 14'h2628;
            14'd 6871: out = 14'h2627;
            14'd 6872: out = 14'h2626;
            14'd 6873: out = 14'h2624;
            14'd 6874: out = 14'h2623;
            14'd 6875: out = 14'h2621;
            14'd 6876: out = 14'h2620;
            14'd 6877: out = 14'h261E;
            14'd 6878: out = 14'h261D;
            14'd 6879: out = 14'h261C;
            14'd 6880: out = 14'h261A;
            14'd 6881: out = 14'h2619;
            14'd 6882: out = 14'h2617;
            14'd 6883: out = 14'h2616;
            14'd 6884: out = 14'h2615;
            14'd 6885: out = 14'h2613;
            14'd 6886: out = 14'h2612;
            14'd 6887: out = 14'h2610;
            14'd 6888: out = 14'h260F;
            14'd 6889: out = 14'h260D;
            14'd 6890: out = 14'h260C;
            14'd 6891: out = 14'h260B;
            14'd 6892: out = 14'h2609;
            14'd 6893: out = 14'h2608;
            14'd 6894: out = 14'h2606;
            14'd 6895: out = 14'h2605;
            14'd 6896: out = 14'h2604;
            14'd 6897: out = 14'h2602;
            14'd 6898: out = 14'h2601;
            14'd 6899: out = 14'h25FF;
            14'd 6900: out = 14'h25FE;
            14'd 6901: out = 14'h25FD;
            14'd 6902: out = 14'h25FB;
            14'd 6903: out = 14'h25FA;
            14'd 6904: out = 14'h25F8;
            14'd 6905: out = 14'h25F7;
            14'd 6906: out = 14'h25F5;
            14'd 6907: out = 14'h25F4;
            14'd 6908: out = 14'h25F3;
            14'd 6909: out = 14'h25F1;
            14'd 6910: out = 14'h25F0;
            14'd 6911: out = 14'h25EE;
            14'd 6912: out = 14'h25ED;
            14'd 6913: out = 14'h25EC;
            14'd 6914: out = 14'h25EA;
            14'd 6915: out = 14'h25E9;
            14'd 6916: out = 14'h25E7;
            14'd 6917: out = 14'h25E6;
            14'd 6918: out = 14'h25E5;
            14'd 6919: out = 14'h25E3;
            14'd 6920: out = 14'h25E2;
            14'd 6921: out = 14'h25E0;
            14'd 6922: out = 14'h25DF;
            14'd 6923: out = 14'h25DE;
            14'd 6924: out = 14'h25DC;
            14'd 6925: out = 14'h25DB;
            14'd 6926: out = 14'h25D9;
            14'd 6927: out = 14'h25D8;
            14'd 6928: out = 14'h25D7;
            14'd 6929: out = 14'h25D5;
            14'd 6930: out = 14'h25D4;
            14'd 6931: out = 14'h25D2;
            14'd 6932: out = 14'h25D1;
            14'd 6933: out = 14'h25D0;
            14'd 6934: out = 14'h25CE;
            14'd 6935: out = 14'h25CD;
            14'd 6936: out = 14'h25CB;
            14'd 6937: out = 14'h25CA;
            14'd 6938: out = 14'h25C9;
            14'd 6939: out = 14'h25C7;
            14'd 6940: out = 14'h25C6;
            14'd 6941: out = 14'h25C4;
            14'd 6942: out = 14'h25C3;
            14'd 6943: out = 14'h25C2;
            14'd 6944: out = 14'h25C0;
            14'd 6945: out = 14'h25BF;
            14'd 6946: out = 14'h25BE;
            14'd 6947: out = 14'h25BC;
            14'd 6948: out = 14'h25BB;
            14'd 6949: out = 14'h25B9;
            14'd 6950: out = 14'h25B8;
            14'd 6951: out = 14'h25B7;
            14'd 6952: out = 14'h25B5;
            14'd 6953: out = 14'h25B4;
            14'd 6954: out = 14'h25B2;
            14'd 6955: out = 14'h25B1;
            14'd 6956: out = 14'h25B0;
            14'd 6957: out = 14'h25AE;
            14'd 6958: out = 14'h25AD;
            14'd 6959: out = 14'h25AB;
            14'd 6960: out = 14'h25AA;
            14'd 6961: out = 14'h25A9;
            14'd 6962: out = 14'h25A7;
            14'd 6963: out = 14'h25A6;
            14'd 6964: out = 14'h25A5;
            14'd 6965: out = 14'h25A3;
            14'd 6966: out = 14'h25A2;
            14'd 6967: out = 14'h25A0;
            14'd 6968: out = 14'h259F;
            14'd 6969: out = 14'h259E;
            14'd 6970: out = 14'h259C;
            14'd 6971: out = 14'h259B;
            14'd 6972: out = 14'h2599;
            14'd 6973: out = 14'h2598;
            14'd 6974: out = 14'h2597;
            14'd 6975: out = 14'h2595;
            14'd 6976: out = 14'h2594;
            14'd 6977: out = 14'h2593;
            14'd 6978: out = 14'h2591;
            14'd 6979: out = 14'h2590;
            14'd 6980: out = 14'h258E;
            14'd 6981: out = 14'h258D;
            14'd 6982: out = 14'h258C;
            14'd 6983: out = 14'h258A;
            14'd 6984: out = 14'h2589;
            14'd 6985: out = 14'h2588;
            14'd 6986: out = 14'h2586;
            14'd 6987: out = 14'h2585;
            14'd 6988: out = 14'h2583;
            14'd 6989: out = 14'h2582;
            14'd 6990: out = 14'h2581;
            14'd 6991: out = 14'h257F;
            14'd 6992: out = 14'h257E;
            14'd 6993: out = 14'h257D;
            14'd 6994: out = 14'h257B;
            14'd 6995: out = 14'h257A;
            14'd 6996: out = 14'h2578;
            14'd 6997: out = 14'h2577;
            14'd 6998: out = 14'h2576;
            14'd 6999: out = 14'h2574;
            14'd 7000: out = 14'h2573;
            14'd 7001: out = 14'h2572;
            14'd 7002: out = 14'h2570;
            14'd 7003: out = 14'h256F;
            14'd 7004: out = 14'h256E;
            14'd 7005: out = 14'h256C;
            14'd 7006: out = 14'h256B;
            14'd 7007: out = 14'h2569;
            14'd 7008: out = 14'h2568;
            14'd 7009: out = 14'h2567;
            14'd 7010: out = 14'h2565;
            14'd 7011: out = 14'h2564;
            14'd 7012: out = 14'h2563;
            14'd 7013: out = 14'h2561;
            14'd 7014: out = 14'h2560;
            14'd 7015: out = 14'h255E;
            14'd 7016: out = 14'h255D;
            14'd 7017: out = 14'h255C;
            14'd 7018: out = 14'h255A;
            14'd 7019: out = 14'h2559;
            14'd 7020: out = 14'h2558;
            14'd 7021: out = 14'h2556;
            14'd 7022: out = 14'h2555;
            14'd 7023: out = 14'h2554;
            14'd 7024: out = 14'h2552;
            14'd 7025: out = 14'h2551;
            14'd 7026: out = 14'h2550;
            14'd 7027: out = 14'h254E;
            14'd 7028: out = 14'h254D;
            14'd 7029: out = 14'h254B;
            14'd 7030: out = 14'h254A;
            14'd 7031: out = 14'h2549;
            14'd 7032: out = 14'h2547;
            14'd 7033: out = 14'h2546;
            14'd 7034: out = 14'h2545;
            14'd 7035: out = 14'h2543;
            14'd 7036: out = 14'h2542;
            14'd 7037: out = 14'h2541;
            14'd 7038: out = 14'h253F;
            14'd 7039: out = 14'h253E;
            14'd 7040: out = 14'h253D;
            14'd 7041: out = 14'h253B;
            14'd 7042: out = 14'h253A;
            14'd 7043: out = 14'h2538;
            14'd 7044: out = 14'h2537;
            14'd 7045: out = 14'h2536;
            14'd 7046: out = 14'h2534;
            14'd 7047: out = 14'h2533;
            14'd 7048: out = 14'h2532;
            14'd 7049: out = 14'h2530;
            14'd 7050: out = 14'h252F;
            14'd 7051: out = 14'h252E;
            14'd 7052: out = 14'h252C;
            14'd 7053: out = 14'h252B;
            14'd 7054: out = 14'h252A;
            14'd 7055: out = 14'h2528;
            14'd 7056: out = 14'h2527;
            14'd 7057: out = 14'h2526;
            14'd 7058: out = 14'h2524;
            14'd 7059: out = 14'h2523;
            14'd 7060: out = 14'h2522;
            14'd 7061: out = 14'h2520;
            14'd 7062: out = 14'h251F;
            14'd 7063: out = 14'h251D;
            14'd 7064: out = 14'h251C;
            14'd 7065: out = 14'h251B;
            14'd 7066: out = 14'h2519;
            14'd 7067: out = 14'h2518;
            14'd 7068: out = 14'h2517;
            14'd 7069: out = 14'h2515;
            14'd 7070: out = 14'h2514;
            14'd 7071: out = 14'h2513;
            14'd 7072: out = 14'h2511;
            14'd 7073: out = 14'h2510;
            14'd 7074: out = 14'h250F;
            14'd 7075: out = 14'h250D;
            14'd 7076: out = 14'h250C;
            14'd 7077: out = 14'h250B;
            14'd 7078: out = 14'h2509;
            14'd 7079: out = 14'h2508;
            14'd 7080: out = 14'h2507;
            14'd 7081: out = 14'h2505;
            14'd 7082: out = 14'h2504;
            14'd 7083: out = 14'h2503;
            14'd 7084: out = 14'h2501;
            14'd 7085: out = 14'h2500;
            14'd 7086: out = 14'h24FF;
            14'd 7087: out = 14'h24FD;
            14'd 7088: out = 14'h24FC;
            14'd 7089: out = 14'h24FB;
            14'd 7090: out = 14'h24F9;
            14'd 7091: out = 14'h24F8;
            14'd 7092: out = 14'h24F7;
            14'd 7093: out = 14'h24F5;
            14'd 7094: out = 14'h24F4;
            14'd 7095: out = 14'h24F3;
            14'd 7096: out = 14'h24F1;
            14'd 7097: out = 14'h24F0;
            14'd 7098: out = 14'h24EF;
            14'd 7099: out = 14'h24ED;
            14'd 7100: out = 14'h24EC;
            14'd 7101: out = 14'h24EB;
            14'd 7102: out = 14'h24E9;
            14'd 7103: out = 14'h24E8;
            14'd 7104: out = 14'h24E7;
            14'd 7105: out = 14'h24E5;
            14'd 7106: out = 14'h24E4;
            14'd 7107: out = 14'h24E3;
            14'd 7108: out = 14'h24E1;
            14'd 7109: out = 14'h24E0;
            14'd 7110: out = 14'h24DF;
            14'd 7111: out = 14'h24DD;
            14'd 7112: out = 14'h24DC;
            14'd 7113: out = 14'h24DB;
            14'd 7114: out = 14'h24D9;
            14'd 7115: out = 14'h24D8;
            14'd 7116: out = 14'h24D7;
            14'd 7117: out = 14'h24D5;
            14'd 7118: out = 14'h24D4;
            14'd 7119: out = 14'h24D3;
            14'd 7120: out = 14'h24D1;
            14'd 7121: out = 14'h24D0;
            14'd 7122: out = 14'h24CF;
            14'd 7123: out = 14'h24CD;
            14'd 7124: out = 14'h24CC;
            14'd 7125: out = 14'h24CB;
            14'd 7126: out = 14'h24C9;
            14'd 7127: out = 14'h24C8;
            14'd 7128: out = 14'h24C7;
            14'd 7129: out = 14'h24C6;
            14'd 7130: out = 14'h24C4;
            14'd 7131: out = 14'h24C3;
            14'd 7132: out = 14'h24C2;
            14'd 7133: out = 14'h24C0;
            14'd 7134: out = 14'h24BF;
            14'd 7135: out = 14'h24BE;
            14'd 7136: out = 14'h24BC;
            14'd 7137: out = 14'h24BB;
            14'd 7138: out = 14'h24BA;
            14'd 7139: out = 14'h24B8;
            14'd 7140: out = 14'h24B7;
            14'd 7141: out = 14'h24B6;
            14'd 7142: out = 14'h24B4;
            14'd 7143: out = 14'h24B3;
            14'd 7144: out = 14'h24B2;
            14'd 7145: out = 14'h24B0;
            14'd 7146: out = 14'h24AF;
            14'd 7147: out = 14'h24AE;
            14'd 7148: out = 14'h24AC;
            14'd 7149: out = 14'h24AB;
            14'd 7150: out = 14'h24AA;
            14'd 7151: out = 14'h24A9;
            14'd 7152: out = 14'h24A7;
            14'd 7153: out = 14'h24A6;
            14'd 7154: out = 14'h24A5;
            14'd 7155: out = 14'h24A3;
            14'd 7156: out = 14'h24A2;
            14'd 7157: out = 14'h24A1;
            14'd 7158: out = 14'h249F;
            14'd 7159: out = 14'h249E;
            14'd 7160: out = 14'h249D;
            14'd 7161: out = 14'h249B;
            14'd 7162: out = 14'h249A;
            14'd 7163: out = 14'h2499;
            14'd 7164: out = 14'h2498;
            14'd 7165: out = 14'h2496;
            14'd 7166: out = 14'h2495;
            14'd 7167: out = 14'h2494;
            14'd 7168: out = 14'h2492;
            14'd 7169: out = 14'h2491;
            14'd 7170: out = 14'h2490;
            14'd 7171: out = 14'h248E;
            14'd 7172: out = 14'h248D;
            14'd 7173: out = 14'h248C;
            14'd 7174: out = 14'h248A;
            14'd 7175: out = 14'h2489;
            14'd 7176: out = 14'h2488;
            14'd 7177: out = 14'h2487;
            14'd 7178: out = 14'h2485;
            14'd 7179: out = 14'h2484;
            14'd 7180: out = 14'h2483;
            14'd 7181: out = 14'h2481;
            14'd 7182: out = 14'h2480;
            14'd 7183: out = 14'h247F;
            14'd 7184: out = 14'h247D;
            14'd 7185: out = 14'h247C;
            14'd 7186: out = 14'h247B;
            14'd 7187: out = 14'h247A;
            14'd 7188: out = 14'h2478;
            14'd 7189: out = 14'h2477;
            14'd 7190: out = 14'h2476;
            14'd 7191: out = 14'h2474;
            14'd 7192: out = 14'h2473;
            14'd 7193: out = 14'h2472;
            14'd 7194: out = 14'h2470;
            14'd 7195: out = 14'h246F;
            14'd 7196: out = 14'h246E;
            14'd 7197: out = 14'h246D;
            14'd 7198: out = 14'h246B;
            14'd 7199: out = 14'h246A;
            14'd 7200: out = 14'h2469;
            14'd 7201: out = 14'h2467;
            14'd 7202: out = 14'h2466;
            14'd 7203: out = 14'h2465;
            14'd 7204: out = 14'h2464;
            14'd 7205: out = 14'h2462;
            14'd 7206: out = 14'h2461;
            14'd 7207: out = 14'h2460;
            14'd 7208: out = 14'h245E;
            14'd 7209: out = 14'h245D;
            14'd 7210: out = 14'h245C;
            14'd 7211: out = 14'h245A;
            14'd 7212: out = 14'h2459;
            14'd 7213: out = 14'h2458;
            14'd 7214: out = 14'h2457;
            14'd 7215: out = 14'h2455;
            14'd 7216: out = 14'h2454;
            14'd 7217: out = 14'h2453;
            14'd 7218: out = 14'h2451;
            14'd 7219: out = 14'h2450;
            14'd 7220: out = 14'h244F;
            14'd 7221: out = 14'h244E;
            14'd 7222: out = 14'h244C;
            14'd 7223: out = 14'h244B;
            14'd 7224: out = 14'h244A;
            14'd 7225: out = 14'h2448;
            14'd 7226: out = 14'h2447;
            14'd 7227: out = 14'h2446;
            14'd 7228: out = 14'h2445;
            14'd 7229: out = 14'h2443;
            14'd 7230: out = 14'h2442;
            14'd 7231: out = 14'h2441;
            14'd 7232: out = 14'h243F;
            14'd 7233: out = 14'h243E;
            14'd 7234: out = 14'h243D;
            14'd 7235: out = 14'h243C;
            14'd 7236: out = 14'h243A;
            14'd 7237: out = 14'h2439;
            14'd 7238: out = 14'h2438;
            14'd 7239: out = 14'h2436;
            14'd 7240: out = 14'h2435;
            14'd 7241: out = 14'h2434;
            14'd 7242: out = 14'h2433;
            14'd 7243: out = 14'h2431;
            14'd 7244: out = 14'h2430;
            14'd 7245: out = 14'h242F;
            14'd 7246: out = 14'h242E;
            14'd 7247: out = 14'h242C;
            14'd 7248: out = 14'h242B;
            14'd 7249: out = 14'h242A;
            14'd 7250: out = 14'h2428;
            14'd 7251: out = 14'h2427;
            14'd 7252: out = 14'h2426;
            14'd 7253: out = 14'h2425;
            14'd 7254: out = 14'h2423;
            14'd 7255: out = 14'h2422;
            14'd 7256: out = 14'h2421;
            14'd 7257: out = 14'h241F;
            14'd 7258: out = 14'h241E;
            14'd 7259: out = 14'h241D;
            14'd 7260: out = 14'h241C;
            14'd 7261: out = 14'h241A;
            14'd 7262: out = 14'h2419;
            14'd 7263: out = 14'h2418;
            14'd 7264: out = 14'h2417;
            14'd 7265: out = 14'h2415;
            14'd 7266: out = 14'h2414;
            14'd 7267: out = 14'h2413;
            14'd 7268: out = 14'h2411;
            14'd 7269: out = 14'h2410;
            14'd 7270: out = 14'h240F;
            14'd 7271: out = 14'h240E;
            14'd 7272: out = 14'h240C;
            14'd 7273: out = 14'h240B;
            14'd 7274: out = 14'h240A;
            14'd 7275: out = 14'h2409;
            14'd 7276: out = 14'h2407;
            14'd 7277: out = 14'h2406;
            14'd 7278: out = 14'h2405;
            14'd 7279: out = 14'h2404;
            14'd 7280: out = 14'h2402;
            14'd 7281: out = 14'h2401;
            14'd 7282: out = 14'h2400;
            14'd 7283: out = 14'h23FE;
            14'd 7284: out = 14'h23FD;
            14'd 7285: out = 14'h23FC;
            14'd 7286: out = 14'h23FB;
            14'd 7287: out = 14'h23F9;
            14'd 7288: out = 14'h23F8;
            14'd 7289: out = 14'h23F7;
            14'd 7290: out = 14'h23F6;
            14'd 7291: out = 14'h23F4;
            14'd 7292: out = 14'h23F3;
            14'd 7293: out = 14'h23F2;
            14'd 7294: out = 14'h23F1;
            14'd 7295: out = 14'h23EF;
            14'd 7296: out = 14'h23EE;
            14'd 7297: out = 14'h23ED;
            14'd 7298: out = 14'h23EC;
            14'd 7299: out = 14'h23EA;
            14'd 7300: out = 14'h23E9;
            14'd 7301: out = 14'h23E8;
            14'd 7302: out = 14'h23E6;
            14'd 7303: out = 14'h23E5;
            14'd 7304: out = 14'h23E4;
            14'd 7305: out = 14'h23E3;
            14'd 7306: out = 14'h23E1;
            14'd 7307: out = 14'h23E0;
            14'd 7308: out = 14'h23DF;
            14'd 7309: out = 14'h23DE;
            14'd 7310: out = 14'h23DC;
            14'd 7311: out = 14'h23DB;
            14'd 7312: out = 14'h23DA;
            14'd 7313: out = 14'h23D9;
            14'd 7314: out = 14'h23D7;
            14'd 7315: out = 14'h23D6;
            14'd 7316: out = 14'h23D5;
            14'd 7317: out = 14'h23D4;
            14'd 7318: out = 14'h23D2;
            14'd 7319: out = 14'h23D1;
            14'd 7320: out = 14'h23D0;
            14'd 7321: out = 14'h23CF;
            14'd 7322: out = 14'h23CD;
            14'd 7323: out = 14'h23CC;
            14'd 7324: out = 14'h23CB;
            14'd 7325: out = 14'h23CA;
            14'd 7326: out = 14'h23C8;
            14'd 7327: out = 14'h23C7;
            14'd 7328: out = 14'h23C6;
            14'd 7329: out = 14'h23C5;
            14'd 7330: out = 14'h23C3;
            14'd 7331: out = 14'h23C2;
            14'd 7332: out = 14'h23C1;
            14'd 7333: out = 14'h23C0;
            14'd 7334: out = 14'h23BE;
            14'd 7335: out = 14'h23BD;
            14'd 7336: out = 14'h23BC;
            14'd 7337: out = 14'h23BB;
            14'd 7338: out = 14'h23B9;
            14'd 7339: out = 14'h23B8;
            14'd 7340: out = 14'h23B7;
            14'd 7341: out = 14'h23B6;
            14'd 7342: out = 14'h23B4;
            14'd 7343: out = 14'h23B3;
            14'd 7344: out = 14'h23B2;
            14'd 7345: out = 14'h23B1;
            14'd 7346: out = 14'h23AF;
            14'd 7347: out = 14'h23AE;
            14'd 7348: out = 14'h23AD;
            14'd 7349: out = 14'h23AC;
            14'd 7350: out = 14'h23AA;
            14'd 7351: out = 14'h23A9;
            14'd 7352: out = 14'h23A8;
            14'd 7353: out = 14'h23A7;
            14'd 7354: out = 14'h23A5;
            14'd 7355: out = 14'h23A4;
            14'd 7356: out = 14'h23A3;
            14'd 7357: out = 14'h23A2;
            14'd 7358: out = 14'h23A1;
            14'd 7359: out = 14'h239F;
            14'd 7360: out = 14'h239E;
            14'd 7361: out = 14'h239D;
            14'd 7362: out = 14'h239C;
            14'd 7363: out = 14'h239A;
            14'd 7364: out = 14'h2399;
            14'd 7365: out = 14'h2398;
            14'd 7366: out = 14'h2397;
            14'd 7367: out = 14'h2395;
            14'd 7368: out = 14'h2394;
            14'd 7369: out = 14'h2393;
            14'd 7370: out = 14'h2392;
            14'd 7371: out = 14'h2390;
            14'd 7372: out = 14'h238F;
            14'd 7373: out = 14'h238E;
            14'd 7374: out = 14'h238D;
            14'd 7375: out = 14'h238C;
            14'd 7376: out = 14'h238A;
            14'd 7377: out = 14'h2389;
            14'd 7378: out = 14'h2388;
            14'd 7379: out = 14'h2387;
            14'd 7380: out = 14'h2385;
            14'd 7381: out = 14'h2384;
            14'd 7382: out = 14'h2383;
            14'd 7383: out = 14'h2382;
            14'd 7384: out = 14'h2380;
            14'd 7385: out = 14'h237F;
            14'd 7386: out = 14'h237E;
            14'd 7387: out = 14'h237D;
            14'd 7388: out = 14'h237B;
            14'd 7389: out = 14'h237A;
            14'd 7390: out = 14'h2379;
            14'd 7391: out = 14'h2378;
            14'd 7392: out = 14'h2377;
            14'd 7393: out = 14'h2375;
            14'd 7394: out = 14'h2374;
            14'd 7395: out = 14'h2373;
            14'd 7396: out = 14'h2372;
            14'd 7397: out = 14'h2370;
            14'd 7398: out = 14'h236F;
            14'd 7399: out = 14'h236E;
            14'd 7400: out = 14'h236D;
            14'd 7401: out = 14'h236C;
            14'd 7402: out = 14'h236A;
            14'd 7403: out = 14'h2369;
            14'd 7404: out = 14'h2368;
            14'd 7405: out = 14'h2367;
            14'd 7406: out = 14'h2365;
            14'd 7407: out = 14'h2364;
            14'd 7408: out = 14'h2363;
            14'd 7409: out = 14'h2362;
            14'd 7410: out = 14'h2361;
            14'd 7411: out = 14'h235F;
            14'd 7412: out = 14'h235E;
            14'd 7413: out = 14'h235D;
            14'd 7414: out = 14'h235C;
            14'd 7415: out = 14'h235A;
            14'd 7416: out = 14'h2359;
            14'd 7417: out = 14'h2358;
            14'd 7418: out = 14'h2357;
            14'd 7419: out = 14'h2356;
            14'd 7420: out = 14'h2354;
            14'd 7421: out = 14'h2353;
            14'd 7422: out = 14'h2352;
            14'd 7423: out = 14'h2351;
            14'd 7424: out = 14'h234F;
            14'd 7425: out = 14'h234E;
            14'd 7426: out = 14'h234D;
            14'd 7427: out = 14'h234C;
            14'd 7428: out = 14'h234B;
            14'd 7429: out = 14'h2349;
            14'd 7430: out = 14'h2348;
            14'd 7431: out = 14'h2347;
            14'd 7432: out = 14'h2346;
            14'd 7433: out = 14'h2345;
            14'd 7434: out = 14'h2343;
            14'd 7435: out = 14'h2342;
            14'd 7436: out = 14'h2341;
            14'd 7437: out = 14'h2340;
            14'd 7438: out = 14'h233E;
            14'd 7439: out = 14'h233D;
            14'd 7440: out = 14'h233C;
            14'd 7441: out = 14'h233B;
            14'd 7442: out = 14'h233A;
            14'd 7443: out = 14'h2338;
            14'd 7444: out = 14'h2337;
            14'd 7445: out = 14'h2336;
            14'd 7446: out = 14'h2335;
            14'd 7447: out = 14'h2334;
            14'd 7448: out = 14'h2332;
            14'd 7449: out = 14'h2331;
            14'd 7450: out = 14'h2330;
            14'd 7451: out = 14'h232F;
            14'd 7452: out = 14'h232D;
            14'd 7453: out = 14'h232C;
            14'd 7454: out = 14'h232B;
            14'd 7455: out = 14'h232A;
            14'd 7456: out = 14'h2329;
            14'd 7457: out = 14'h2327;
            14'd 7458: out = 14'h2326;
            14'd 7459: out = 14'h2325;
            14'd 7460: out = 14'h2324;
            14'd 7461: out = 14'h2323;
            14'd 7462: out = 14'h2321;
            14'd 7463: out = 14'h2320;
            14'd 7464: out = 14'h231F;
            14'd 7465: out = 14'h231E;
            14'd 7466: out = 14'h231D;
            14'd 7467: out = 14'h231B;
            14'd 7468: out = 14'h231A;
            14'd 7469: out = 14'h2319;
            14'd 7470: out = 14'h2318;
            14'd 7471: out = 14'h2317;
            14'd 7472: out = 14'h2315;
            14'd 7473: out = 14'h2314;
            14'd 7474: out = 14'h2313;
            14'd 7475: out = 14'h2312;
            14'd 7476: out = 14'h2311;
            14'd 7477: out = 14'h230F;
            14'd 7478: out = 14'h230E;
            14'd 7479: out = 14'h230D;
            14'd 7480: out = 14'h230C;
            14'd 7481: out = 14'h230B;
            14'd 7482: out = 14'h2309;
            14'd 7483: out = 14'h2308;
            14'd 7484: out = 14'h2307;
            14'd 7485: out = 14'h2306;
            14'd 7486: out = 14'h2305;
            14'd 7487: out = 14'h2303;
            14'd 7488: out = 14'h2302;
            14'd 7489: out = 14'h2301;
            14'd 7490: out = 14'h2300;
            14'd 7491: out = 14'h22FF;
            14'd 7492: out = 14'h22FD;
            14'd 7493: out = 14'h22FC;
            14'd 7494: out = 14'h22FB;
            14'd 7495: out = 14'h22FA;
            14'd 7496: out = 14'h22F9;
            14'd 7497: out = 14'h22F7;
            14'd 7498: out = 14'h22F6;
            14'd 7499: out = 14'h22F5;
            14'd 7500: out = 14'h22F4;
            14'd 7501: out = 14'h22F3;
            14'd 7502: out = 14'h22F1;
            14'd 7503: out = 14'h22F0;
            14'd 7504: out = 14'h22EF;
            14'd 7505: out = 14'h22EE;
            14'd 7506: out = 14'h22ED;
            14'd 7507: out = 14'h22EC;
            14'd 7508: out = 14'h22EA;
            14'd 7509: out = 14'h22E9;
            14'd 7510: out = 14'h22E8;
            14'd 7511: out = 14'h22E7;
            14'd 7512: out = 14'h22E6;
            14'd 7513: out = 14'h22E4;
            14'd 7514: out = 14'h22E3;
            14'd 7515: out = 14'h22E2;
            14'd 7516: out = 14'h22E1;
            14'd 7517: out = 14'h22E0;
            14'd 7518: out = 14'h22DE;
            14'd 7519: out = 14'h22DD;
            14'd 7520: out = 14'h22DC;
            14'd 7521: out = 14'h22DB;
            14'd 7522: out = 14'h22DA;
            14'd 7523: out = 14'h22D8;
            14'd 7524: out = 14'h22D7;
            14'd 7525: out = 14'h22D6;
            14'd 7526: out = 14'h22D5;
            14'd 7527: out = 14'h22D4;
            14'd 7528: out = 14'h22D3;
            14'd 7529: out = 14'h22D1;
            14'd 7530: out = 14'h22D0;
            14'd 7531: out = 14'h22CF;
            14'd 7532: out = 14'h22CE;
            14'd 7533: out = 14'h22CD;
            14'd 7534: out = 14'h22CB;
            14'd 7535: out = 14'h22CA;
            14'd 7536: out = 14'h22C9;
            14'd 7537: out = 14'h22C8;
            14'd 7538: out = 14'h22C7;
            14'd 7539: out = 14'h22C6;
            14'd 7540: out = 14'h22C4;
            14'd 7541: out = 14'h22C3;
            14'd 7542: out = 14'h22C2;
            14'd 7543: out = 14'h22C1;
            14'd 7544: out = 14'h22C0;
            14'd 7545: out = 14'h22BE;
            14'd 7546: out = 14'h22BD;
            14'd 7547: out = 14'h22BC;
            14'd 7548: out = 14'h22BB;
            14'd 7549: out = 14'h22BA;
            14'd 7550: out = 14'h22B9;
            14'd 7551: out = 14'h22B7;
            14'd 7552: out = 14'h22B6;
            14'd 7553: out = 14'h22B5;
            14'd 7554: out = 14'h22B4;
            14'd 7555: out = 14'h22B3;
            14'd 7556: out = 14'h22B2;
            14'd 7557: out = 14'h22B0;
            14'd 7558: out = 14'h22AF;
            14'd 7559: out = 14'h22AE;
            14'd 7560: out = 14'h22AD;
            14'd 7561: out = 14'h22AC;
            14'd 7562: out = 14'h22AA;
            14'd 7563: out = 14'h22A9;
            14'd 7564: out = 14'h22A8;
            14'd 7565: out = 14'h22A7;
            14'd 7566: out = 14'h22A6;
            14'd 7567: out = 14'h22A5;
            14'd 7568: out = 14'h22A3;
            14'd 7569: out = 14'h22A2;
            14'd 7570: out = 14'h22A1;
            14'd 7571: out = 14'h22A0;
            14'd 7572: out = 14'h229F;
            14'd 7573: out = 14'h229E;
            14'd 7574: out = 14'h229C;
            14'd 7575: out = 14'h229B;
            14'd 7576: out = 14'h229A;
            14'd 7577: out = 14'h2299;
            14'd 7578: out = 14'h2298;
            14'd 7579: out = 14'h2297;
            14'd 7580: out = 14'h2295;
            14'd 7581: out = 14'h2294;
            14'd 7582: out = 14'h2293;
            14'd 7583: out = 14'h2292;
            14'd 7584: out = 14'h2291;
            14'd 7585: out = 14'h2290;
            14'd 7586: out = 14'h228E;
            14'd 7587: out = 14'h228D;
            14'd 7588: out = 14'h228C;
            14'd 7589: out = 14'h228B;
            14'd 7590: out = 14'h228A;
            14'd 7591: out = 14'h2289;
            14'd 7592: out = 14'h2287;
            14'd 7593: out = 14'h2286;
            14'd 7594: out = 14'h2285;
            14'd 7595: out = 14'h2284;
            14'd 7596: out = 14'h2283;
            14'd 7597: out = 14'h2282;
            14'd 7598: out = 14'h2280;
            14'd 7599: out = 14'h227F;
            14'd 7600: out = 14'h227E;
            14'd 7601: out = 14'h227D;
            14'd 7602: out = 14'h227C;
            14'd 7603: out = 14'h227B;
            14'd 7604: out = 14'h2279;
            14'd 7605: out = 14'h2278;
            14'd 7606: out = 14'h2277;
            14'd 7607: out = 14'h2276;
            14'd 7608: out = 14'h2275;
            14'd 7609: out = 14'h2274;
            14'd 7610: out = 14'h2273;
            14'd 7611: out = 14'h2271;
            14'd 7612: out = 14'h2270;
            14'd 7613: out = 14'h226F;
            14'd 7614: out = 14'h226E;
            14'd 7615: out = 14'h226D;
            14'd 7616: out = 14'h226C;
            14'd 7617: out = 14'h226A;
            14'd 7618: out = 14'h2269;
            14'd 7619: out = 14'h2268;
            14'd 7620: out = 14'h2267;
            14'd 7621: out = 14'h2266;
            14'd 7622: out = 14'h2265;
            14'd 7623: out = 14'h2263;
            14'd 7624: out = 14'h2262;
            14'd 7625: out = 14'h2261;
            14'd 7626: out = 14'h2260;
            14'd 7627: out = 14'h225F;
            14'd 7628: out = 14'h225E;
            14'd 7629: out = 14'h225D;
            14'd 7630: out = 14'h225B;
            14'd 7631: out = 14'h225A;
            14'd 7632: out = 14'h2259;
            14'd 7633: out = 14'h2258;
            14'd 7634: out = 14'h2257;
            14'd 7635: out = 14'h2256;
            14'd 7636: out = 14'h2254;
            14'd 7637: out = 14'h2253;
            14'd 7638: out = 14'h2252;
            14'd 7639: out = 14'h2251;
            14'd 7640: out = 14'h2250;
            14'd 7641: out = 14'h224F;
            14'd 7642: out = 14'h224E;
            14'd 7643: out = 14'h224C;
            14'd 7644: out = 14'h224B;
            14'd 7645: out = 14'h224A;
            14'd 7646: out = 14'h2249;
            14'd 7647: out = 14'h2248;
            14'd 7648: out = 14'h2247;
            14'd 7649: out = 14'h2246;
            14'd 7650: out = 14'h2244;
            14'd 7651: out = 14'h2243;
            14'd 7652: out = 14'h2242;
            14'd 7653: out = 14'h2241;
            14'd 7654: out = 14'h2240;
            14'd 7655: out = 14'h223F;
            14'd 7656: out = 14'h223E;
            14'd 7657: out = 14'h223C;
            14'd 7658: out = 14'h223B;
            14'd 7659: out = 14'h223A;
            14'd 7660: out = 14'h2239;
            14'd 7661: out = 14'h2238;
            14'd 7662: out = 14'h2237;
            14'd 7663: out = 14'h2236;
            14'd 7664: out = 14'h2234;
            14'd 7665: out = 14'h2233;
            14'd 7666: out = 14'h2232;
            14'd 7667: out = 14'h2231;
            14'd 7668: out = 14'h2230;
            14'd 7669: out = 14'h222F;
            14'd 7670: out = 14'h222E;
            14'd 7671: out = 14'h222C;
            14'd 7672: out = 14'h222B;
            14'd 7673: out = 14'h222A;
            14'd 7674: out = 14'h2229;
            14'd 7675: out = 14'h2228;
            14'd 7676: out = 14'h2227;
            14'd 7677: out = 14'h2226;
            14'd 7678: out = 14'h2224;
            14'd 7679: out = 14'h2223;
            14'd 7680: out = 14'h2222;
            14'd 7681: out = 14'h2221;
            14'd 7682: out = 14'h2220;
            14'd 7683: out = 14'h221F;
            14'd 7684: out = 14'h221E;
            14'd 7685: out = 14'h221C;
            14'd 7686: out = 14'h221B;
            14'd 7687: out = 14'h221A;
            14'd 7688: out = 14'h2219;
            14'd 7689: out = 14'h2218;
            14'd 7690: out = 14'h2217;
            14'd 7691: out = 14'h2216;
            14'd 7692: out = 14'h2215;
            14'd 7693: out = 14'h2213;
            14'd 7694: out = 14'h2212;
            14'd 7695: out = 14'h2211;
            14'd 7696: out = 14'h2210;
            14'd 7697: out = 14'h220F;
            14'd 7698: out = 14'h220E;
            14'd 7699: out = 14'h220D;
            14'd 7700: out = 14'h220B;
            14'd 7701: out = 14'h220A;
            14'd 7702: out = 14'h2209;
            14'd 7703: out = 14'h2208;
            14'd 7704: out = 14'h2207;
            14'd 7705: out = 14'h2206;
            14'd 7706: out = 14'h2205;
            14'd 7707: out = 14'h2204;
            14'd 7708: out = 14'h2202;
            14'd 7709: out = 14'h2201;
            14'd 7710: out = 14'h2200;
            14'd 7711: out = 14'h21FF;
            14'd 7712: out = 14'h21FE;
            14'd 7713: out = 14'h21FD;
            14'd 7714: out = 14'h21FC;
            14'd 7715: out = 14'h21FA;
            14'd 7716: out = 14'h21F9;
            14'd 7717: out = 14'h21F8;
            14'd 7718: out = 14'h21F7;
            14'd 7719: out = 14'h21F6;
            14'd 7720: out = 14'h21F5;
            14'd 7721: out = 14'h21F4;
            14'd 7722: out = 14'h21F3;
            14'd 7723: out = 14'h21F1;
            14'd 7724: out = 14'h21F0;
            14'd 7725: out = 14'h21EF;
            14'd 7726: out = 14'h21EE;
            14'd 7727: out = 14'h21ED;
            14'd 7728: out = 14'h21EC;
            14'd 7729: out = 14'h21EB;
            14'd 7730: out = 14'h21EA;
            14'd 7731: out = 14'h21E8;
            14'd 7732: out = 14'h21E7;
            14'd 7733: out = 14'h21E6;
            14'd 7734: out = 14'h21E5;
            14'd 7735: out = 14'h21E4;
            14'd 7736: out = 14'h21E3;
            14'd 7737: out = 14'h21E2;
            14'd 7738: out = 14'h21E1;
            14'd 7739: out = 14'h21E0;
            14'd 7740: out = 14'h21DE;
            14'd 7741: out = 14'h21DD;
            14'd 7742: out = 14'h21DC;
            14'd 7743: out = 14'h21DB;
            14'd 7744: out = 14'h21DA;
            14'd 7745: out = 14'h21D9;
            14'd 7746: out = 14'h21D8;
            14'd 7747: out = 14'h21D7;
            14'd 7748: out = 14'h21D5;
            14'd 7749: out = 14'h21D4;
            14'd 7750: out = 14'h21D3;
            14'd 7751: out = 14'h21D2;
            14'd 7752: out = 14'h21D1;
            14'd 7753: out = 14'h21D0;
            14'd 7754: out = 14'h21CF;
            14'd 7755: out = 14'h21CE;
            14'd 7756: out = 14'h21CD;
            14'd 7757: out = 14'h21CB;
            14'd 7758: out = 14'h21CA;
            14'd 7759: out = 14'h21C9;
            14'd 7760: out = 14'h21C8;
            14'd 7761: out = 14'h21C7;
            14'd 7762: out = 14'h21C6;
            14'd 7763: out = 14'h21C5;
            14'd 7764: out = 14'h21C4;
            14'd 7765: out = 14'h21C2;
            14'd 7766: out = 14'h21C1;
            14'd 7767: out = 14'h21C0;
            14'd 7768: out = 14'h21BF;
            14'd 7769: out = 14'h21BE;
            14'd 7770: out = 14'h21BD;
            14'd 7771: out = 14'h21BC;
            14'd 7772: out = 14'h21BB;
            14'd 7773: out = 14'h21BA;
            14'd 7774: out = 14'h21B8;
            14'd 7775: out = 14'h21B7;
            14'd 7776: out = 14'h21B6;
            14'd 7777: out = 14'h21B5;
            14'd 7778: out = 14'h21B4;
            14'd 7779: out = 14'h21B3;
            14'd 7780: out = 14'h21B2;
            14'd 7781: out = 14'h21B1;
            14'd 7782: out = 14'h21B0;
            14'd 7783: out = 14'h21AE;
            14'd 7784: out = 14'h21AD;
            14'd 7785: out = 14'h21AC;
            14'd 7786: out = 14'h21AB;
            14'd 7787: out = 14'h21AA;
            14'd 7788: out = 14'h21A9;
            14'd 7789: out = 14'h21A8;
            14'd 7790: out = 14'h21A7;
            14'd 7791: out = 14'h21A6;
            14'd 7792: out = 14'h21A5;
            14'd 7793: out = 14'h21A3;
            14'd 7794: out = 14'h21A2;
            14'd 7795: out = 14'h21A1;
            14'd 7796: out = 14'h21A0;
            14'd 7797: out = 14'h219F;
            14'd 7798: out = 14'h219E;
            14'd 7799: out = 14'h219D;
            14'd 7800: out = 14'h219C;
            14'd 7801: out = 14'h219B;
            14'd 7802: out = 14'h2199;
            14'd 7803: out = 14'h2198;
            14'd 7804: out = 14'h2197;
            14'd 7805: out = 14'h2196;
            14'd 7806: out = 14'h2195;
            14'd 7807: out = 14'h2194;
            14'd 7808: out = 14'h2193;
            14'd 7809: out = 14'h2192;
            14'd 7810: out = 14'h2191;
            14'd 7811: out = 14'h2190;
            14'd 7812: out = 14'h218E;
            14'd 7813: out = 14'h218D;
            14'd 7814: out = 14'h218C;
            14'd 7815: out = 14'h218B;
            14'd 7816: out = 14'h218A;
            14'd 7817: out = 14'h2189;
            14'd 7818: out = 14'h2188;
            14'd 7819: out = 14'h2187;
            14'd 7820: out = 14'h2186;
            14'd 7821: out = 14'h2185;
            14'd 7822: out = 14'h2184;
            14'd 7823: out = 14'h2182;
            14'd 7824: out = 14'h2181;
            14'd 7825: out = 14'h2180;
            14'd 7826: out = 14'h217F;
            14'd 7827: out = 14'h217E;
            14'd 7828: out = 14'h217D;
            14'd 7829: out = 14'h217C;
            14'd 7830: out = 14'h217B;
            14'd 7831: out = 14'h217A;
            14'd 7832: out = 14'h2179;
            14'd 7833: out = 14'h2177;
            14'd 7834: out = 14'h2176;
            14'd 7835: out = 14'h2175;
            14'd 7836: out = 14'h2174;
            14'd 7837: out = 14'h2173;
            14'd 7838: out = 14'h2172;
            14'd 7839: out = 14'h2171;
            14'd 7840: out = 14'h2170;
            14'd 7841: out = 14'h216F;
            14'd 7842: out = 14'h216E;
            14'd 7843: out = 14'h216D;
            14'd 7844: out = 14'h216B;
            14'd 7845: out = 14'h216A;
            14'd 7846: out = 14'h2169;
            14'd 7847: out = 14'h2168;
            14'd 7848: out = 14'h2167;
            14'd 7849: out = 14'h2166;
            14'd 7850: out = 14'h2165;
            14'd 7851: out = 14'h2164;
            14'd 7852: out = 14'h2163;
            14'd 7853: out = 14'h2162;
            14'd 7854: out = 14'h2161;
            14'd 7855: out = 14'h215F;
            14'd 7856: out = 14'h215E;
            14'd 7857: out = 14'h215D;
            14'd 7858: out = 14'h215C;
            14'd 7859: out = 14'h215B;
            14'd 7860: out = 14'h215A;
            14'd 7861: out = 14'h2159;
            14'd 7862: out = 14'h2158;
            14'd 7863: out = 14'h2157;
            14'd 7864: out = 14'h2156;
            14'd 7865: out = 14'h2155;
            14'd 7866: out = 14'h2154;
            14'd 7867: out = 14'h2152;
            14'd 7868: out = 14'h2151;
            14'd 7869: out = 14'h2150;
            14'd 7870: out = 14'h214F;
            14'd 7871: out = 14'h214E;
            14'd 7872: out = 14'h214D;
            14'd 7873: out = 14'h214C;
            14'd 7874: out = 14'h214B;
            14'd 7875: out = 14'h214A;
            14'd 7876: out = 14'h2149;
            14'd 7877: out = 14'h2148;
            14'd 7878: out = 14'h2147;
            14'd 7879: out = 14'h2145;
            14'd 7880: out = 14'h2144;
            14'd 7881: out = 14'h2143;
            14'd 7882: out = 14'h2142;
            14'd 7883: out = 14'h2141;
            14'd 7884: out = 14'h2140;
            14'd 7885: out = 14'h213F;
            14'd 7886: out = 14'h213E;
            14'd 7887: out = 14'h213D;
            14'd 7888: out = 14'h213C;
            14'd 7889: out = 14'h213B;
            14'd 7890: out = 14'h213A;
            14'd 7891: out = 14'h2138;
            14'd 7892: out = 14'h2137;
            14'd 7893: out = 14'h2136;
            14'd 7894: out = 14'h2135;
            14'd 7895: out = 14'h2134;
            14'd 7896: out = 14'h2133;
            14'd 7897: out = 14'h2132;
            14'd 7898: out = 14'h2131;
            14'd 7899: out = 14'h2130;
            14'd 7900: out = 14'h212F;
            14'd 7901: out = 14'h212E;
            14'd 7902: out = 14'h212D;
            14'd 7903: out = 14'h212C;
            14'd 7904: out = 14'h212A;
            14'd 7905: out = 14'h2129;
            14'd 7906: out = 14'h2128;
            14'd 7907: out = 14'h2127;
            14'd 7908: out = 14'h2126;
            14'd 7909: out = 14'h2125;
            14'd 7910: out = 14'h2124;
            14'd 7911: out = 14'h2123;
            14'd 7912: out = 14'h2122;
            14'd 7913: out = 14'h2121;
            14'd 7914: out = 14'h2120;
            14'd 7915: out = 14'h211F;
            14'd 7916: out = 14'h211E;
            14'd 7917: out = 14'h211D;
            14'd 7918: out = 14'h211B;
            14'd 7919: out = 14'h211A;
            14'd 7920: out = 14'h2119;
            14'd 7921: out = 14'h2118;
            14'd 7922: out = 14'h2117;
            14'd 7923: out = 14'h2116;
            14'd 7924: out = 14'h2115;
            14'd 7925: out = 14'h2114;
            14'd 7926: out = 14'h2113;
            14'd 7927: out = 14'h2112;
            14'd 7928: out = 14'h2111;
            14'd 7929: out = 14'h2110;
            14'd 7930: out = 14'h210F;
            14'd 7931: out = 14'h210E;
            14'd 7932: out = 14'h210D;
            14'd 7933: out = 14'h210B;
            14'd 7934: out = 14'h210A;
            14'd 7935: out = 14'h2109;
            14'd 7936: out = 14'h2108;
            14'd 7937: out = 14'h2107;
            14'd 7938: out = 14'h2106;
            14'd 7939: out = 14'h2105;
            14'd 7940: out = 14'h2104;
            14'd 7941: out = 14'h2103;
            14'd 7942: out = 14'h2102;
            14'd 7943: out = 14'h2101;
            14'd 7944: out = 14'h2100;
            14'd 7945: out = 14'h20FF;
            14'd 7946: out = 14'h20FE;
            14'd 7947: out = 14'h20FD;
            14'd 7948: out = 14'h20FB;
            14'd 7949: out = 14'h20FA;
            14'd 7950: out = 14'h20F9;
            14'd 7951: out = 14'h20F8;
            14'd 7952: out = 14'h20F7;
            14'd 7953: out = 14'h20F6;
            14'd 7954: out = 14'h20F5;
            14'd 7955: out = 14'h20F4;
            14'd 7956: out = 14'h20F3;
            14'd 7957: out = 14'h20F2;
            14'd 7958: out = 14'h20F1;
            14'd 7959: out = 14'h20F0;
            14'd 7960: out = 14'h20EF;
            14'd 7961: out = 14'h20EE;
            14'd 7962: out = 14'h20ED;
            14'd 7963: out = 14'h20EC;
            14'd 7964: out = 14'h20EB;
            14'd 7965: out = 14'h20E9;
            14'd 7966: out = 14'h20E8;
            14'd 7967: out = 14'h20E7;
            14'd 7968: out = 14'h20E6;
            14'd 7969: out = 14'h20E5;
            14'd 7970: out = 14'h20E4;
            14'd 7971: out = 14'h20E3;
            14'd 7972: out = 14'h20E2;
            14'd 7973: out = 14'h20E1;
            14'd 7974: out = 14'h20E0;
            14'd 7975: out = 14'h20DF;
            14'd 7976: out = 14'h20DE;
            14'd 7977: out = 14'h20DD;
            14'd 7978: out = 14'h20DC;
            14'd 7979: out = 14'h20DB;
            14'd 7980: out = 14'h20DA;
            14'd 7981: out = 14'h20D9;
            14'd 7982: out = 14'h20D8;
            14'd 7983: out = 14'h20D6;
            14'd 7984: out = 14'h20D5;
            14'd 7985: out = 14'h20D4;
            14'd 7986: out = 14'h20D3;
            14'd 7987: out = 14'h20D2;
            14'd 7988: out = 14'h20D1;
            14'd 7989: out = 14'h20D0;
            14'd 7990: out = 14'h20CF;
            14'd 7991: out = 14'h20CE;
            14'd 7992: out = 14'h20CD;
            14'd 7993: out = 14'h20CC;
            14'd 7994: out = 14'h20CB;
            14'd 7995: out = 14'h20CA;
            14'd 7996: out = 14'h20C9;
            14'd 7997: out = 14'h20C8;
            14'd 7998: out = 14'h20C7;
            14'd 7999: out = 14'h20C6;
            14'd 8000: out = 14'h20C5;
            14'd 8001: out = 14'h20C4;
            14'd 8002: out = 14'h20C3;
            14'd 8003: out = 14'h20C1;
            14'd 8004: out = 14'h20C0;
            14'd 8005: out = 14'h20BF;
            14'd 8006: out = 14'h20BE;
            14'd 8007: out = 14'h20BD;
            14'd 8008: out = 14'h20BC;
            14'd 8009: out = 14'h20BB;
            14'd 8010: out = 14'h20BA;
            14'd 8011: out = 14'h20B9;
            14'd 8012: out = 14'h20B8;
            14'd 8013: out = 14'h20B7;
            14'd 8014: out = 14'h20B6;
            14'd 8015: out = 14'h20B5;
            14'd 8016: out = 14'h20B4;
            14'd 8017: out = 14'h20B3;
            14'd 8018: out = 14'h20B2;
            14'd 8019: out = 14'h20B1;
            14'd 8020: out = 14'h20B0;
            14'd 8021: out = 14'h20AF;
            14'd 8022: out = 14'h20AE;
            14'd 8023: out = 14'h20AD;
            14'd 8024: out = 14'h20AC;
            14'd 8025: out = 14'h20AA;
            14'd 8026: out = 14'h20A9;
            14'd 8027: out = 14'h20A8;
            14'd 8028: out = 14'h20A7;
            14'd 8029: out = 14'h20A6;
            14'd 8030: out = 14'h20A5;
            14'd 8031: out = 14'h20A4;
            14'd 8032: out = 14'h20A3;
            14'd 8033: out = 14'h20A2;
            14'd 8034: out = 14'h20A1;
            14'd 8035: out = 14'h20A0;
            14'd 8036: out = 14'h209F;
            14'd 8037: out = 14'h209E;
            14'd 8038: out = 14'h209D;
            14'd 8039: out = 14'h209C;
            14'd 8040: out = 14'h209B;
            14'd 8041: out = 14'h209A;
            14'd 8042: out = 14'h2099;
            14'd 8043: out = 14'h2098;
            14'd 8044: out = 14'h2097;
            14'd 8045: out = 14'h2096;
            14'd 8046: out = 14'h2095;
            14'd 8047: out = 14'h2094;
            14'd 8048: out = 14'h2093;
            14'd 8049: out = 14'h2092;
            14'd 8050: out = 14'h2091;
            14'd 8051: out = 14'h208F;
            14'd 8052: out = 14'h208E;
            14'd 8053: out = 14'h208D;
            14'd 8054: out = 14'h208C;
            14'd 8055: out = 14'h208B;
            14'd 8056: out = 14'h208A;
            14'd 8057: out = 14'h2089;
            14'd 8058: out = 14'h2088;
            14'd 8059: out = 14'h2087;
            14'd 8060: out = 14'h2086;
            14'd 8061: out = 14'h2085;
            14'd 8062: out = 14'h2084;
            14'd 8063: out = 14'h2083;
            14'd 8064: out = 14'h2082;
            14'd 8065: out = 14'h2081;
            14'd 8066: out = 14'h2080;
            14'd 8067: out = 14'h207F;
            14'd 8068: out = 14'h207E;
            14'd 8069: out = 14'h207D;
            14'd 8070: out = 14'h207C;
            14'd 8071: out = 14'h207B;
            14'd 8072: out = 14'h207A;
            14'd 8073: out = 14'h2079;
            14'd 8074: out = 14'h2078;
            14'd 8075: out = 14'h2077;
            14'd 8076: out = 14'h2076;
            14'd 8077: out = 14'h2075;
            14'd 8078: out = 14'h2074;
            14'd 8079: out = 14'h2073;
            14'd 8080: out = 14'h2072;
            14'd 8081: out = 14'h2071;
            14'd 8082: out = 14'h206F;
            14'd 8083: out = 14'h206E;
            14'd 8084: out = 14'h206D;
            14'd 8085: out = 14'h206C;
            14'd 8086: out = 14'h206B;
            14'd 8087: out = 14'h206A;
            14'd 8088: out = 14'h2069;
            14'd 8089: out = 14'h2068;
            14'd 8090: out = 14'h2067;
            14'd 8091: out = 14'h2066;
            14'd 8092: out = 14'h2065;
            14'd 8093: out = 14'h2064;
            14'd 8094: out = 14'h2063;
            14'd 8095: out = 14'h2062;
            14'd 8096: out = 14'h2061;
            14'd 8097: out = 14'h2060;
            14'd 8098: out = 14'h205F;
            14'd 8099: out = 14'h205E;
            14'd 8100: out = 14'h205D;
            14'd 8101: out = 14'h205C;
            14'd 8102: out = 14'h205B;
            14'd 8103: out = 14'h205A;
            14'd 8104: out = 14'h2059;
            14'd 8105: out = 14'h2058;
            14'd 8106: out = 14'h2057;
            14'd 8107: out = 14'h2056;
            14'd 8108: out = 14'h2055;
            14'd 8109: out = 14'h2054;
            14'd 8110: out = 14'h2053;
            14'd 8111: out = 14'h2052;
            14'd 8112: out = 14'h2051;
            14'd 8113: out = 14'h2050;
            14'd 8114: out = 14'h204F;
            14'd 8115: out = 14'h204E;
            14'd 8116: out = 14'h204D;
            14'd 8117: out = 14'h204C;
            14'd 8118: out = 14'h204B;
            14'd 8119: out = 14'h204A;
            14'd 8120: out = 14'h2049;
            14'd 8121: out = 14'h2048;
            14'd 8122: out = 14'h2047;
            14'd 8123: out = 14'h2046;
            14'd 8124: out = 14'h2045;
            14'd 8125: out = 14'h2044;
            14'd 8126: out = 14'h2043;
            14'd 8127: out = 14'h2042;
            14'd 8128: out = 14'h2041;
            14'd 8129: out = 14'h203F;
            14'd 8130: out = 14'h203E;
            14'd 8131: out = 14'h203D;
            14'd 8132: out = 14'h203C;
            14'd 8133: out = 14'h203B;
            14'd 8134: out = 14'h203A;
            14'd 8135: out = 14'h2039;
            14'd 8136: out = 14'h2038;
            14'd 8137: out = 14'h2037;
            14'd 8138: out = 14'h2036;
            14'd 8139: out = 14'h2035;
            14'd 8140: out = 14'h2034;
            14'd 8141: out = 14'h2033;
            14'd 8142: out = 14'h2032;
            14'd 8143: out = 14'h2031;
            14'd 8144: out = 14'h2030;
            14'd 8145: out = 14'h202F;
            14'd 8146: out = 14'h202E;
            14'd 8147: out = 14'h202D;
            14'd 8148: out = 14'h202C;
            14'd 8149: out = 14'h202B;
            14'd 8150: out = 14'h202A;
            14'd 8151: out = 14'h2029;
            14'd 8152: out = 14'h2028;
            14'd 8153: out = 14'h2027;
            14'd 8154: out = 14'h2026;
            14'd 8155: out = 14'h2025;
            14'd 8156: out = 14'h2024;
            14'd 8157: out = 14'h2023;
            14'd 8158: out = 14'h2022;
            14'd 8159: out = 14'h2021;
            14'd 8160: out = 14'h2020;
            14'd 8161: out = 14'h201F;
            14'd 8162: out = 14'h201E;
            14'd 8163: out = 14'h201D;
            14'd 8164: out = 14'h201C;
            14'd 8165: out = 14'h201B;
            14'd 8166: out = 14'h201A;
            14'd 8167: out = 14'h2019;
            14'd 8168: out = 14'h2018;
            14'd 8169: out = 14'h2017;
            14'd 8170: out = 14'h2016;
            14'd 8171: out = 14'h2015;
            14'd 8172: out = 14'h2014;
            14'd 8173: out = 14'h2013;
            14'd 8174: out = 14'h2012;
            14'd 8175: out = 14'h2011;
            14'd 8176: out = 14'h2010;
            14'd 8177: out = 14'h200F;
            14'd 8178: out = 14'h200E;
            14'd 8179: out = 14'h200D;
            14'd 8180: out = 14'h200C;
            14'd 8181: out = 14'h200B;
            14'd 8182: out = 14'h200A;
            14'd 8183: out = 14'h2009;
            14'd 8184: out = 14'h2008;
            14'd 8185: out = 14'h2007;
            14'd 8186: out = 14'h2006;
            14'd 8187: out = 14'h2005;
            14'd 8188: out = 14'h2004;
            14'd 8189: out = 14'h2003;
            14'd 8190: out = 14'h2002;
            14'd 8191: out = 14'h2001;
            14'd 8192: out = 14'h2000;
            14'd 8193: out = 14'h1FFF;
            14'd 8194: out = 14'h1FFE;
            14'd 8195: out = 14'h1FFD;
            14'd 8196: out = 14'h1FFC;
            14'd 8197: out = 14'h1FFB;
            14'd 8198: out = 14'h1FFA;
            14'd 8199: out = 14'h1FF9;
            14'd 8200: out = 14'h1FF8;
            14'd 8201: out = 14'h1FF7;
            14'd 8202: out = 14'h1FF6;
            14'd 8203: out = 14'h1FF5;
            14'd 8204: out = 14'h1FF4;
            14'd 8205: out = 14'h1FF3;
            14'd 8206: out = 14'h1FF2;
            14'd 8207: out = 14'h1FF1;
            14'd 8208: out = 14'h1FF0;
            14'd 8209: out = 14'h1FEF;
            14'd 8210: out = 14'h1FEE;
            14'd 8211: out = 14'h1FED;
            14'd 8212: out = 14'h1FEC;
            14'd 8213: out = 14'h1FEB;
            14'd 8214: out = 14'h1FEA;
            14'd 8215: out = 14'h1FE9;
            14'd 8216: out = 14'h1FE8;
            14'd 8217: out = 14'h1FE7;
            14'd 8218: out = 14'h1FE6;
            14'd 8219: out = 14'h1FE5;
            14'd 8220: out = 14'h1FE4;
            14'd 8221: out = 14'h1FE3;
            14'd 8222: out = 14'h1FE2;
            14'd 8223: out = 14'h1FE1;
            14'd 8224: out = 14'h1FE0;
            14'd 8225: out = 14'h1FDF;
            14'd 8226: out = 14'h1FDE;
            14'd 8227: out = 14'h1FDD;
            14'd 8228: out = 14'h1FDC;
            14'd 8229: out = 14'h1FDB;
            14'd 8230: out = 14'h1FDA;
            14'd 8231: out = 14'h1FD9;
            14'd 8232: out = 14'h1FD8;
            14'd 8233: out = 14'h1FD7;
            14'd 8234: out = 14'h1FD6;
            14'd 8235: out = 14'h1FD5;
            14'd 8236: out = 14'h1FD4;
            14'd 8237: out = 14'h1FD3;
            14'd 8238: out = 14'h1FD2;
            14'd 8239: out = 14'h1FD1;
            14'd 8240: out = 14'h1FD0;
            14'd 8241: out = 14'h1FCF;
            14'd 8242: out = 14'h1FCE;
            14'd 8243: out = 14'h1FCD;
            14'd 8244: out = 14'h1FCC;
            14'd 8245: out = 14'h1FCB;
            14'd 8246: out = 14'h1FCA;
            14'd 8247: out = 14'h1FC9;
            14'd 8248: out = 14'h1FC8;
            14'd 8249: out = 14'h1FC7;
            14'd 8250: out = 14'h1FC6;
            14'd 8251: out = 14'h1FC5;
            14'd 8252: out = 14'h1FC4;
            14'd 8253: out = 14'h1FC3;
            14'd 8254: out = 14'h1FC2;
            14'd 8255: out = 14'h1FC1;
            14'd 8256: out = 14'h1FC0;
            14'd 8257: out = 14'h1FC0;
            14'd 8258: out = 14'h1FBF;
            14'd 8259: out = 14'h1FBE;
            14'd 8260: out = 14'h1FBD;
            14'd 8261: out = 14'h1FBC;
            14'd 8262: out = 14'h1FBB;
            14'd 8263: out = 14'h1FBA;
            14'd 8264: out = 14'h1FB9;
            14'd 8265: out = 14'h1FB8;
            14'd 8266: out = 14'h1FB7;
            14'd 8267: out = 14'h1FB6;
            14'd 8268: out = 14'h1FB5;
            14'd 8269: out = 14'h1FB4;
            14'd 8270: out = 14'h1FB3;
            14'd 8271: out = 14'h1FB2;
            14'd 8272: out = 14'h1FB1;
            14'd 8273: out = 14'h1FB0;
            14'd 8274: out = 14'h1FAF;
            14'd 8275: out = 14'h1FAE;
            14'd 8276: out = 14'h1FAD;
            14'd 8277: out = 14'h1FAC;
            14'd 8278: out = 14'h1FAB;
            14'd 8279: out = 14'h1FAA;
            14'd 8280: out = 14'h1FA9;
            14'd 8281: out = 14'h1FA8;
            14'd 8282: out = 14'h1FA7;
            14'd 8283: out = 14'h1FA6;
            14'd 8284: out = 14'h1FA5;
            14'd 8285: out = 14'h1FA4;
            14'd 8286: out = 14'h1FA3;
            14'd 8287: out = 14'h1FA2;
            14'd 8288: out = 14'h1FA1;
            14'd 8289: out = 14'h1FA0;
            14'd 8290: out = 14'h1F9F;
            14'd 8291: out = 14'h1F9E;
            14'd 8292: out = 14'h1F9D;
            14'd 8293: out = 14'h1F9C;
            14'd 8294: out = 14'h1F9B;
            14'd 8295: out = 14'h1F9A;
            14'd 8296: out = 14'h1F99;
            14'd 8297: out = 14'h1F98;
            14'd 8298: out = 14'h1F97;
            14'd 8299: out = 14'h1F96;
            14'd 8300: out = 14'h1F95;
            14'd 8301: out = 14'h1F94;
            14'd 8302: out = 14'h1F93;
            14'd 8303: out = 14'h1F92;
            14'd 8304: out = 14'h1F92;
            14'd 8305: out = 14'h1F91;
            14'd 8306: out = 14'h1F90;
            14'd 8307: out = 14'h1F8F;
            14'd 8308: out = 14'h1F8E;
            14'd 8309: out = 14'h1F8D;
            14'd 8310: out = 14'h1F8C;
            14'd 8311: out = 14'h1F8B;
            14'd 8312: out = 14'h1F8A;
            14'd 8313: out = 14'h1F89;
            14'd 8314: out = 14'h1F88;
            14'd 8315: out = 14'h1F87;
            14'd 8316: out = 14'h1F86;
            14'd 8317: out = 14'h1F85;
            14'd 8318: out = 14'h1F84;
            14'd 8319: out = 14'h1F83;
            14'd 8320: out = 14'h1F82;
            14'd 8321: out = 14'h1F81;
            14'd 8322: out = 14'h1F80;
            14'd 8323: out = 14'h1F7F;
            14'd 8324: out = 14'h1F7E;
            14'd 8325: out = 14'h1F7D;
            14'd 8326: out = 14'h1F7C;
            14'd 8327: out = 14'h1F7B;
            14'd 8328: out = 14'h1F7A;
            14'd 8329: out = 14'h1F79;
            14'd 8330: out = 14'h1F78;
            14'd 8331: out = 14'h1F77;
            14'd 8332: out = 14'h1F76;
            14'd 8333: out = 14'h1F75;
            14'd 8334: out = 14'h1F74;
            14'd 8335: out = 14'h1F73;
            14'd 8336: out = 14'h1F72;
            14'd 8337: out = 14'h1F72;
            14'd 8338: out = 14'h1F71;
            14'd 8339: out = 14'h1F70;
            14'd 8340: out = 14'h1F6F;
            14'd 8341: out = 14'h1F6E;
            14'd 8342: out = 14'h1F6D;
            14'd 8343: out = 14'h1F6C;
            14'd 8344: out = 14'h1F6B;
            14'd 8345: out = 14'h1F6A;
            14'd 8346: out = 14'h1F69;
            14'd 8347: out = 14'h1F68;
            14'd 8348: out = 14'h1F67;
            14'd 8349: out = 14'h1F66;
            14'd 8350: out = 14'h1F65;
            14'd 8351: out = 14'h1F64;
            14'd 8352: out = 14'h1F63;
            14'd 8353: out = 14'h1F62;
            14'd 8354: out = 14'h1F61;
            14'd 8355: out = 14'h1F60;
            14'd 8356: out = 14'h1F5F;
            14'd 8357: out = 14'h1F5E;
            14'd 8358: out = 14'h1F5D;
            14'd 8359: out = 14'h1F5C;
            14'd 8360: out = 14'h1F5B;
            14'd 8361: out = 14'h1F5A;
            14'd 8362: out = 14'h1F59;
            14'd 8363: out = 14'h1F58;
            14'd 8364: out = 14'h1F58;
            14'd 8365: out = 14'h1F57;
            14'd 8366: out = 14'h1F56;
            14'd 8367: out = 14'h1F55;
            14'd 8368: out = 14'h1F54;
            14'd 8369: out = 14'h1F53;
            14'd 8370: out = 14'h1F52;
            14'd 8371: out = 14'h1F51;
            14'd 8372: out = 14'h1F50;
            14'd 8373: out = 14'h1F4F;
            14'd 8374: out = 14'h1F4E;
            14'd 8375: out = 14'h1F4D;
            14'd 8376: out = 14'h1F4C;
            14'd 8377: out = 14'h1F4B;
            14'd 8378: out = 14'h1F4A;
            14'd 8379: out = 14'h1F49;
            14'd 8380: out = 14'h1F48;
            14'd 8381: out = 14'h1F47;
            14'd 8382: out = 14'h1F46;
            14'd 8383: out = 14'h1F45;
            14'd 8384: out = 14'h1F44;
            14'd 8385: out = 14'h1F43;
            14'd 8386: out = 14'h1F42;
            14'd 8387: out = 14'h1F42;
            14'd 8388: out = 14'h1F41;
            14'd 8389: out = 14'h1F40;
            14'd 8390: out = 14'h1F3F;
            14'd 8391: out = 14'h1F3E;
            14'd 8392: out = 14'h1F3D;
            14'd 8393: out = 14'h1F3C;
            14'd 8394: out = 14'h1F3B;
            14'd 8395: out = 14'h1F3A;
            14'd 8396: out = 14'h1F39;
            14'd 8397: out = 14'h1F38;
            14'd 8398: out = 14'h1F37;
            14'd 8399: out = 14'h1F36;
            14'd 8400: out = 14'h1F35;
            14'd 8401: out = 14'h1F34;
            14'd 8402: out = 14'h1F33;
            14'd 8403: out = 14'h1F32;
            14'd 8404: out = 14'h1F31;
            14'd 8405: out = 14'h1F30;
            14'd 8406: out = 14'h1F2F;
            14'd 8407: out = 14'h1F2E;
            14'd 8408: out = 14'h1F2E;
            14'd 8409: out = 14'h1F2D;
            14'd 8410: out = 14'h1F2C;
            14'd 8411: out = 14'h1F2B;
            14'd 8412: out = 14'h1F2A;
            14'd 8413: out = 14'h1F29;
            14'd 8414: out = 14'h1F28;
            14'd 8415: out = 14'h1F27;
            14'd 8416: out = 14'h1F26;
            14'd 8417: out = 14'h1F25;
            14'd 8418: out = 14'h1F24;
            14'd 8419: out = 14'h1F23;
            14'd 8420: out = 14'h1F22;
            14'd 8421: out = 14'h1F21;
            14'd 8422: out = 14'h1F20;
            14'd 8423: out = 14'h1F1F;
            14'd 8424: out = 14'h1F1E;
            14'd 8425: out = 14'h1F1D;
            14'd 8426: out = 14'h1F1C;
            14'd 8427: out = 14'h1F1C;
            14'd 8428: out = 14'h1F1B;
            14'd 8429: out = 14'h1F1A;
            14'd 8430: out = 14'h1F19;
            14'd 8431: out = 14'h1F18;
            14'd 8432: out = 14'h1F17;
            14'd 8433: out = 14'h1F16;
            14'd 8434: out = 14'h1F15;
            14'd 8435: out = 14'h1F14;
            14'd 8436: out = 14'h1F13;
            14'd 8437: out = 14'h1F12;
            14'd 8438: out = 14'h1F11;
            14'd 8439: out = 14'h1F10;
            14'd 8440: out = 14'h1F0F;
            14'd 8441: out = 14'h1F0E;
            14'd 8442: out = 14'h1F0D;
            14'd 8443: out = 14'h1F0C;
            14'd 8444: out = 14'h1F0C;
            14'd 8445: out = 14'h1F0B;
            14'd 8446: out = 14'h1F0A;
            14'd 8447: out = 14'h1F09;
            14'd 8448: out = 14'h1F08;
            14'd 8449: out = 14'h1F07;
            14'd 8450: out = 14'h1F06;
            14'd 8451: out = 14'h1F05;
            14'd 8452: out = 14'h1F04;
            14'd 8453: out = 14'h1F03;
            14'd 8454: out = 14'h1F02;
            14'd 8455: out = 14'h1F01;
            14'd 8456: out = 14'h1F00;
            14'd 8457: out = 14'h1EFF;
            14'd 8458: out = 14'h1EFE;
            14'd 8459: out = 14'h1EFD;
            14'd 8460: out = 14'h1EFC;
            14'd 8461: out = 14'h1EFC;
            14'd 8462: out = 14'h1EFB;
            14'd 8463: out = 14'h1EFA;
            14'd 8464: out = 14'h1EF9;
            14'd 8465: out = 14'h1EF8;
            14'd 8466: out = 14'h1EF7;
            14'd 8467: out = 14'h1EF6;
            14'd 8468: out = 14'h1EF5;
            14'd 8469: out = 14'h1EF4;
            14'd 8470: out = 14'h1EF3;
            14'd 8471: out = 14'h1EF2;
            14'd 8472: out = 14'h1EF1;
            14'd 8473: out = 14'h1EF0;
            14'd 8474: out = 14'h1EEF;
            14'd 8475: out = 14'h1EEE;
            14'd 8476: out = 14'h1EEE;
            14'd 8477: out = 14'h1EED;
            14'd 8478: out = 14'h1EEC;
            14'd 8479: out = 14'h1EEB;
            14'd 8480: out = 14'h1EEA;
            14'd 8481: out = 14'h1EE9;
            14'd 8482: out = 14'h1EE8;
            14'd 8483: out = 14'h1EE7;
            14'd 8484: out = 14'h1EE6;
            14'd 8485: out = 14'h1EE5;
            14'd 8486: out = 14'h1EE4;
            14'd 8487: out = 14'h1EE3;
            14'd 8488: out = 14'h1EE2;
            14'd 8489: out = 14'h1EE1;
            14'd 8490: out = 14'h1EE0;
            14'd 8491: out = 14'h1EE0;
            14'd 8492: out = 14'h1EDF;
            14'd 8493: out = 14'h1EDE;
            14'd 8494: out = 14'h1EDD;
            14'd 8495: out = 14'h1EDC;
            14'd 8496: out = 14'h1EDB;
            14'd 8497: out = 14'h1EDA;
            14'd 8498: out = 14'h1ED9;
            14'd 8499: out = 14'h1ED8;
            14'd 8500: out = 14'h1ED7;
            14'd 8501: out = 14'h1ED6;
            14'd 8502: out = 14'h1ED5;
            14'd 8503: out = 14'h1ED4;
            14'd 8504: out = 14'h1ED3;
            14'd 8505: out = 14'h1ED3;
            14'd 8506: out = 14'h1ED2;
            14'd 8507: out = 14'h1ED1;
            14'd 8508: out = 14'h1ED0;
            14'd 8509: out = 14'h1ECF;
            14'd 8510: out = 14'h1ECE;
            14'd 8511: out = 14'h1ECD;
            14'd 8512: out = 14'h1ECC;
            14'd 8513: out = 14'h1ECB;
            14'd 8514: out = 14'h1ECA;
            14'd 8515: out = 14'h1EC9;
            14'd 8516: out = 14'h1EC8;
            14'd 8517: out = 14'h1EC7;
            14'd 8518: out = 14'h1EC6;
            14'd 8519: out = 14'h1EC6;
            14'd 8520: out = 14'h1EC5;
            14'd 8521: out = 14'h1EC4;
            14'd 8522: out = 14'h1EC3;
            14'd 8523: out = 14'h1EC2;
            14'd 8524: out = 14'h1EC1;
            14'd 8525: out = 14'h1EC0;
            14'd 8526: out = 14'h1EBF;
            14'd 8527: out = 14'h1EBE;
            14'd 8528: out = 14'h1EBD;
            14'd 8529: out = 14'h1EBC;
            14'd 8530: out = 14'h1EBB;
            14'd 8531: out = 14'h1EBA;
            14'd 8532: out = 14'h1EBA;
            14'd 8533: out = 14'h1EB9;
            14'd 8534: out = 14'h1EB8;
            14'd 8535: out = 14'h1EB7;
            14'd 8536: out = 14'h1EB6;
            14'd 8537: out = 14'h1EB5;
            14'd 8538: out = 14'h1EB4;
            14'd 8539: out = 14'h1EB3;
            14'd 8540: out = 14'h1EB2;
            14'd 8541: out = 14'h1EB1;
            14'd 8542: out = 14'h1EB0;
            14'd 8543: out = 14'h1EAF;
            14'd 8544: out = 14'h1EAF;
            14'd 8545: out = 14'h1EAE;
            14'd 8546: out = 14'h1EAD;
            14'd 8547: out = 14'h1EAC;
            14'd 8548: out = 14'h1EAB;
            14'd 8549: out = 14'h1EAA;
            14'd 8550: out = 14'h1EA9;
            14'd 8551: out = 14'h1EA8;
            14'd 8552: out = 14'h1EA7;
            14'd 8553: out = 14'h1EA6;
            14'd 8554: out = 14'h1EA5;
            14'd 8555: out = 14'h1EA4;
            14'd 8556: out = 14'h1EA3;
            14'd 8557: out = 14'h1EA3;
            14'd 8558: out = 14'h1EA2;
            14'd 8559: out = 14'h1EA1;
            14'd 8560: out = 14'h1EA0;
            14'd 8561: out = 14'h1E9F;
            14'd 8562: out = 14'h1E9E;
            14'd 8563: out = 14'h1E9D;
            14'd 8564: out = 14'h1E9C;
            14'd 8565: out = 14'h1E9B;
            14'd 8566: out = 14'h1E9A;
            14'd 8567: out = 14'h1E99;
            14'd 8568: out = 14'h1E99;
            14'd 8569: out = 14'h1E98;
            14'd 8570: out = 14'h1E97;
            14'd 8571: out = 14'h1E96;
            14'd 8572: out = 14'h1E95;
            14'd 8573: out = 14'h1E94;
            14'd 8574: out = 14'h1E93;
            14'd 8575: out = 14'h1E92;
            14'd 8576: out = 14'h1E91;
            14'd 8577: out = 14'h1E90;
            14'd 8578: out = 14'h1E8F;
            14'd 8579: out = 14'h1E8E;
            14'd 8580: out = 14'h1E8E;
            14'd 8581: out = 14'h1E8D;
            14'd 8582: out = 14'h1E8C;
            14'd 8583: out = 14'h1E8B;
            14'd 8584: out = 14'h1E8A;
            14'd 8585: out = 14'h1E89;
            14'd 8586: out = 14'h1E88;
            14'd 8587: out = 14'h1E87;
            14'd 8588: out = 14'h1E86;
            14'd 8589: out = 14'h1E85;
            14'd 8590: out = 14'h1E84;
            14'd 8591: out = 14'h1E84;
            14'd 8592: out = 14'h1E83;
            14'd 8593: out = 14'h1E82;
            14'd 8594: out = 14'h1E81;
            14'd 8595: out = 14'h1E80;
            14'd 8596: out = 14'h1E7F;
            14'd 8597: out = 14'h1E7E;
            14'd 8598: out = 14'h1E7D;
            14'd 8599: out = 14'h1E7C;
            14'd 8600: out = 14'h1E7B;
            14'd 8601: out = 14'h1E7A;
            14'd 8602: out = 14'h1E7A;
            14'd 8603: out = 14'h1E79;
            14'd 8604: out = 14'h1E78;
            14'd 8605: out = 14'h1E77;
            14'd 8606: out = 14'h1E76;
            14'd 8607: out = 14'h1E75;
            14'd 8608: out = 14'h1E74;
            14'd 8609: out = 14'h1E73;
            14'd 8610: out = 14'h1E72;
            14'd 8611: out = 14'h1E71;
            14'd 8612: out = 14'h1E70;
            14'd 8613: out = 14'h1E70;
            14'd 8614: out = 14'h1E6F;
            14'd 8615: out = 14'h1E6E;
            14'd 8616: out = 14'h1E6D;
            14'd 8617: out = 14'h1E6C;
            14'd 8618: out = 14'h1E6B;
            14'd 8619: out = 14'h1E6A;
            14'd 8620: out = 14'h1E69;
            14'd 8621: out = 14'h1E68;
            14'd 8622: out = 14'h1E67;
            14'd 8623: out = 14'h1E67;
            14'd 8624: out = 14'h1E66;
            14'd 8625: out = 14'h1E65;
            14'd 8626: out = 14'h1E64;
            14'd 8627: out = 14'h1E63;
            14'd 8628: out = 14'h1E62;
            14'd 8629: out = 14'h1E61;
            14'd 8630: out = 14'h1E60;
            14'd 8631: out = 14'h1E5F;
            14'd 8632: out = 14'h1E5E;
            14'd 8633: out = 14'h1E5E;
            14'd 8634: out = 14'h1E5D;
            14'd 8635: out = 14'h1E5C;
            14'd 8636: out = 14'h1E5B;
            14'd 8637: out = 14'h1E5A;
            14'd 8638: out = 14'h1E59;
            14'd 8639: out = 14'h1E58;
            14'd 8640: out = 14'h1E57;
            14'd 8641: out = 14'h1E56;
            14'd 8642: out = 14'h1E55;
            14'd 8643: out = 14'h1E55;
            14'd 8644: out = 14'h1E54;
            14'd 8645: out = 14'h1E53;
            14'd 8646: out = 14'h1E52;
            14'd 8647: out = 14'h1E51;
            14'd 8648: out = 14'h1E50;
            14'd 8649: out = 14'h1E4F;
            14'd 8650: out = 14'h1E4E;
            14'd 8651: out = 14'h1E4D;
            14'd 8652: out = 14'h1E4C;
            14'd 8653: out = 14'h1E4C;
            14'd 8654: out = 14'h1E4B;
            14'd 8655: out = 14'h1E4A;
            14'd 8656: out = 14'h1E49;
            14'd 8657: out = 14'h1E48;
            14'd 8658: out = 14'h1E47;
            14'd 8659: out = 14'h1E46;
            14'd 8660: out = 14'h1E45;
            14'd 8661: out = 14'h1E44;
            14'd 8662: out = 14'h1E44;
            14'd 8663: out = 14'h1E43;
            14'd 8664: out = 14'h1E42;
            14'd 8665: out = 14'h1E41;
            14'd 8666: out = 14'h1E40;
            14'd 8667: out = 14'h1E3F;
            14'd 8668: out = 14'h1E3E;
            14'd 8669: out = 14'h1E3D;
            14'd 8670: out = 14'h1E3C;
            14'd 8671: out = 14'h1E3B;
            14'd 8672: out = 14'h1E3B;
            14'd 8673: out = 14'h1E3A;
            14'd 8674: out = 14'h1E39;
            14'd 8675: out = 14'h1E38;
            14'd 8676: out = 14'h1E37;
            14'd 8677: out = 14'h1E36;
            14'd 8678: out = 14'h1E35;
            14'd 8679: out = 14'h1E34;
            14'd 8680: out = 14'h1E33;
            14'd 8681: out = 14'h1E33;
            14'd 8682: out = 14'h1E32;
            14'd 8683: out = 14'h1E31;
            14'd 8684: out = 14'h1E30;
            14'd 8685: out = 14'h1E2F;
            14'd 8686: out = 14'h1E2E;
            14'd 8687: out = 14'h1E2D;
            14'd 8688: out = 14'h1E2C;
            14'd 8689: out = 14'h1E2B;
            14'd 8690: out = 14'h1E2B;
            14'd 8691: out = 14'h1E2A;
            14'd 8692: out = 14'h1E29;
            14'd 8693: out = 14'h1E28;
            14'd 8694: out = 14'h1E27;
            14'd 8695: out = 14'h1E26;
            14'd 8696: out = 14'h1E25;
            14'd 8697: out = 14'h1E24;
            14'd 8698: out = 14'h1E23;
            14'd 8699: out = 14'h1E23;
            14'd 8700: out = 14'h1E22;
            14'd 8701: out = 14'h1E21;
            14'd 8702: out = 14'h1E20;
            14'd 8703: out = 14'h1E1F;
            14'd 8704: out = 14'h1E1E;
            14'd 8705: out = 14'h1E1D;
            14'd 8706: out = 14'h1E1C;
            14'd 8707: out = 14'h1E1B;
            14'd 8708: out = 14'h1E1B;
            14'd 8709: out = 14'h1E1A;
            14'd 8710: out = 14'h1E19;
            14'd 8711: out = 14'h1E18;
            14'd 8712: out = 14'h1E17;
            14'd 8713: out = 14'h1E16;
            14'd 8714: out = 14'h1E15;
            14'd 8715: out = 14'h1E14;
            14'd 8716: out = 14'h1E14;
            14'd 8717: out = 14'h1E13;
            14'd 8718: out = 14'h1E12;
            14'd 8719: out = 14'h1E11;
            14'd 8720: out = 14'h1E10;
            14'd 8721: out = 14'h1E0F;
            14'd 8722: out = 14'h1E0E;
            14'd 8723: out = 14'h1E0D;
            14'd 8724: out = 14'h1E0C;
            14'd 8725: out = 14'h1E0C;
            14'd 8726: out = 14'h1E0B;
            14'd 8727: out = 14'h1E0A;
            14'd 8728: out = 14'h1E09;
            14'd 8729: out = 14'h1E08;
            14'd 8730: out = 14'h1E07;
            14'd 8731: out = 14'h1E06;
            14'd 8732: out = 14'h1E05;
            14'd 8733: out = 14'h1E05;
            14'd 8734: out = 14'h1E04;
            14'd 8735: out = 14'h1E03;
            14'd 8736: out = 14'h1E02;
            14'd 8737: out = 14'h1E01;
            14'd 8738: out = 14'h1E00;
            14'd 8739: out = 14'h1DFF;
            14'd 8740: out = 14'h1DFE;
            14'd 8741: out = 14'h1DFD;
            14'd 8742: out = 14'h1DFD;
            14'd 8743: out = 14'h1DFC;
            14'd 8744: out = 14'h1DFB;
            14'd 8745: out = 14'h1DFA;
            14'd 8746: out = 14'h1DF9;
            14'd 8747: out = 14'h1DF8;
            14'd 8748: out = 14'h1DF7;
            14'd 8749: out = 14'h1DF6;
            14'd 8750: out = 14'h1DF6;
            14'd 8751: out = 14'h1DF5;
            14'd 8752: out = 14'h1DF4;
            14'd 8753: out = 14'h1DF3;
            14'd 8754: out = 14'h1DF2;
            14'd 8755: out = 14'h1DF1;
            14'd 8756: out = 14'h1DF0;
            14'd 8757: out = 14'h1DEF;
            14'd 8758: out = 14'h1DEF;
            14'd 8759: out = 14'h1DEE;
            14'd 8760: out = 14'h1DED;
            14'd 8761: out = 14'h1DEC;
            14'd 8762: out = 14'h1DEB;
            14'd 8763: out = 14'h1DEA;
            14'd 8764: out = 14'h1DE9;
            14'd 8765: out = 14'h1DE8;
            14'd 8766: out = 14'h1DE8;
            14'd 8767: out = 14'h1DE7;
            14'd 8768: out = 14'h1DE6;
            14'd 8769: out = 14'h1DE5;
            14'd 8770: out = 14'h1DE4;
            14'd 8771: out = 14'h1DE3;
            14'd 8772: out = 14'h1DE2;
            14'd 8773: out = 14'h1DE1;
            14'd 8774: out = 14'h1DE1;
            14'd 8775: out = 14'h1DE0;
            14'd 8776: out = 14'h1DDF;
            14'd 8777: out = 14'h1DDE;
            14'd 8778: out = 14'h1DDD;
            14'd 8779: out = 14'h1DDC;
            14'd 8780: out = 14'h1DDB;
            14'd 8781: out = 14'h1DDB;
            14'd 8782: out = 14'h1DDA;
            14'd 8783: out = 14'h1DD9;
            14'd 8784: out = 14'h1DD8;
            14'd 8785: out = 14'h1DD7;
            14'd 8786: out = 14'h1DD6;
            14'd 8787: out = 14'h1DD5;
            14'd 8788: out = 14'h1DD4;
            14'd 8789: out = 14'h1DD4;
            14'd 8790: out = 14'h1DD3;
            14'd 8791: out = 14'h1DD2;
            14'd 8792: out = 14'h1DD1;
            14'd 8793: out = 14'h1DD0;
            14'd 8794: out = 14'h1DCF;
            14'd 8795: out = 14'h1DCE;
            14'd 8796: out = 14'h1DCD;
            14'd 8797: out = 14'h1DCD;
            14'd 8798: out = 14'h1DCC;
            14'd 8799: out = 14'h1DCB;
            14'd 8800: out = 14'h1DCA;
            14'd 8801: out = 14'h1DC9;
            14'd 8802: out = 14'h1DC8;
            14'd 8803: out = 14'h1DC7;
            14'd 8804: out = 14'h1DC7;
            14'd 8805: out = 14'h1DC6;
            14'd 8806: out = 14'h1DC5;
            14'd 8807: out = 14'h1DC4;
            14'd 8808: out = 14'h1DC3;
            14'd 8809: out = 14'h1DC2;
            14'd 8810: out = 14'h1DC1;
            14'd 8811: out = 14'h1DC0;
            14'd 8812: out = 14'h1DC0;
            14'd 8813: out = 14'h1DBF;
            14'd 8814: out = 14'h1DBE;
            14'd 8815: out = 14'h1DBD;
            14'd 8816: out = 14'h1DBC;
            14'd 8817: out = 14'h1DBB;
            14'd 8818: out = 14'h1DBA;
            14'd 8819: out = 14'h1DBA;
            14'd 8820: out = 14'h1DB9;
            14'd 8821: out = 14'h1DB8;
            14'd 8822: out = 14'h1DB7;
            14'd 8823: out = 14'h1DB6;
            14'd 8824: out = 14'h1DB5;
            14'd 8825: out = 14'h1DB4;
            14'd 8826: out = 14'h1DB4;
            14'd 8827: out = 14'h1DB3;
            14'd 8828: out = 14'h1DB2;
            14'd 8829: out = 14'h1DB1;
            14'd 8830: out = 14'h1DB0;
            14'd 8831: out = 14'h1DAF;
            14'd 8832: out = 14'h1DAE;
            14'd 8833: out = 14'h1DAE;
            14'd 8834: out = 14'h1DAD;
            14'd 8835: out = 14'h1DAC;
            14'd 8836: out = 14'h1DAB;
            14'd 8837: out = 14'h1DAA;
            14'd 8838: out = 14'h1DA9;
            14'd 8839: out = 14'h1DA8;
            14'd 8840: out = 14'h1DA8;
            14'd 8841: out = 14'h1DA7;
            14'd 8842: out = 14'h1DA6;
            14'd 8843: out = 14'h1DA5;
            14'd 8844: out = 14'h1DA4;
            14'd 8845: out = 14'h1DA3;
            14'd 8846: out = 14'h1DA2;
            14'd 8847: out = 14'h1DA1;
            14'd 8848: out = 14'h1DA1;
            14'd 8849: out = 14'h1DA0;
            14'd 8850: out = 14'h1D9F;
            14'd 8851: out = 14'h1D9E;
            14'd 8852: out = 14'h1D9D;
            14'd 8853: out = 14'h1D9C;
            14'd 8854: out = 14'h1D9B;
            14'd 8855: out = 14'h1D9B;
            14'd 8856: out = 14'h1D9A;
            14'd 8857: out = 14'h1D99;
            14'd 8858: out = 14'h1D98;
            14'd 8859: out = 14'h1D97;
            14'd 8860: out = 14'h1D96;
            14'd 8861: out = 14'h1D96;
            14'd 8862: out = 14'h1D95;
            14'd 8863: out = 14'h1D94;
            14'd 8864: out = 14'h1D93;
            14'd 8865: out = 14'h1D92;
            14'd 8866: out = 14'h1D91;
            14'd 8867: out = 14'h1D90;
            14'd 8868: out = 14'h1D90;
            14'd 8869: out = 14'h1D8F;
            14'd 8870: out = 14'h1D8E;
            14'd 8871: out = 14'h1D8D;
            14'd 8872: out = 14'h1D8C;
            14'd 8873: out = 14'h1D8B;
            14'd 8874: out = 14'h1D8A;
            14'd 8875: out = 14'h1D8A;
            14'd 8876: out = 14'h1D89;
            14'd 8877: out = 14'h1D88;
            14'd 8878: out = 14'h1D87;
            14'd 8879: out = 14'h1D86;
            14'd 8880: out = 14'h1D85;
            14'd 8881: out = 14'h1D84;
            14'd 8882: out = 14'h1D84;
            14'd 8883: out = 14'h1D83;
            14'd 8884: out = 14'h1D82;
            14'd 8885: out = 14'h1D81;
            14'd 8886: out = 14'h1D80;
            14'd 8887: out = 14'h1D7F;
            14'd 8888: out = 14'h1D7F;
            14'd 8889: out = 14'h1D7E;
            14'd 8890: out = 14'h1D7D;
            14'd 8891: out = 14'h1D7C;
            14'd 8892: out = 14'h1D7B;
            14'd 8893: out = 14'h1D7A;
            14'd 8894: out = 14'h1D79;
            14'd 8895: out = 14'h1D79;
            14'd 8896: out = 14'h1D78;
            14'd 8897: out = 14'h1D77;
            14'd 8898: out = 14'h1D76;
            14'd 8899: out = 14'h1D75;
            14'd 8900: out = 14'h1D74;
            14'd 8901: out = 14'h1D73;
            14'd 8902: out = 14'h1D73;
            14'd 8903: out = 14'h1D72;
            14'd 8904: out = 14'h1D71;
            14'd 8905: out = 14'h1D70;
            14'd 8906: out = 14'h1D6F;
            14'd 8907: out = 14'h1D6E;
            14'd 8908: out = 14'h1D6E;
            14'd 8909: out = 14'h1D6D;
            14'd 8910: out = 14'h1D6C;
            14'd 8911: out = 14'h1D6B;
            14'd 8912: out = 14'h1D6A;
            14'd 8913: out = 14'h1D69;
            14'd 8914: out = 14'h1D68;
            14'd 8915: out = 14'h1D68;
            14'd 8916: out = 14'h1D67;
            14'd 8917: out = 14'h1D66;
            14'd 8918: out = 14'h1D65;
            14'd 8919: out = 14'h1D64;
            14'd 8920: out = 14'h1D63;
            14'd 8921: out = 14'h1D63;
            14'd 8922: out = 14'h1D62;
            14'd 8923: out = 14'h1D61;
            14'd 8924: out = 14'h1D60;
            14'd 8925: out = 14'h1D5F;
            14'd 8926: out = 14'h1D5E;
            14'd 8927: out = 14'h1D5E;
            14'd 8928: out = 14'h1D5D;
            14'd 8929: out = 14'h1D5C;
            14'd 8930: out = 14'h1D5B;
            14'd 8931: out = 14'h1D5A;
            14'd 8932: out = 14'h1D59;
            14'd 8933: out = 14'h1D58;
            14'd 8934: out = 14'h1D58;
            14'd 8935: out = 14'h1D57;
            14'd 8936: out = 14'h1D56;
            14'd 8937: out = 14'h1D55;
            14'd 8938: out = 14'h1D54;
            14'd 8939: out = 14'h1D53;
            14'd 8940: out = 14'h1D53;
            14'd 8941: out = 14'h1D52;
            14'd 8942: out = 14'h1D51;
            14'd 8943: out = 14'h1D50;
            14'd 8944: out = 14'h1D4F;
            14'd 8945: out = 14'h1D4E;
            14'd 8946: out = 14'h1D4E;
            14'd 8947: out = 14'h1D4D;
            14'd 8948: out = 14'h1D4C;
            14'd 8949: out = 14'h1D4B;
            14'd 8950: out = 14'h1D4A;
            14'd 8951: out = 14'h1D49;
            14'd 8952: out = 14'h1D49;
            14'd 8953: out = 14'h1D48;
            14'd 8954: out = 14'h1D47;
            14'd 8955: out = 14'h1D46;
            14'd 8956: out = 14'h1D45;
            14'd 8957: out = 14'h1D44;
            14'd 8958: out = 14'h1D44;
            14'd 8959: out = 14'h1D43;
            14'd 8960: out = 14'h1D42;
            14'd 8961: out = 14'h1D41;
            14'd 8962: out = 14'h1D40;
            14'd 8963: out = 14'h1D3F;
            14'd 8964: out = 14'h1D3E;
            14'd 8965: out = 14'h1D3E;
            14'd 8966: out = 14'h1D3D;
            14'd 8967: out = 14'h1D3C;
            14'd 8968: out = 14'h1D3B;
            14'd 8969: out = 14'h1D3A;
            14'd 8970: out = 14'h1D39;
            14'd 8971: out = 14'h1D39;
            14'd 8972: out = 14'h1D38;
            14'd 8973: out = 14'h1D37;
            14'd 8974: out = 14'h1D36;
            14'd 8975: out = 14'h1D35;
            14'd 8976: out = 14'h1D34;
            14'd 8977: out = 14'h1D34;
            14'd 8978: out = 14'h1D33;
            14'd 8979: out = 14'h1D32;
            14'd 8980: out = 14'h1D31;
            14'd 8981: out = 14'h1D30;
            14'd 8982: out = 14'h1D2F;
            14'd 8983: out = 14'h1D2F;
            14'd 8984: out = 14'h1D2E;
            14'd 8985: out = 14'h1D2D;
            14'd 8986: out = 14'h1D2C;
            14'd 8987: out = 14'h1D2B;
            14'd 8988: out = 14'h1D2A;
            14'd 8989: out = 14'h1D2A;
            14'd 8990: out = 14'h1D29;
            14'd 8991: out = 14'h1D28;
            14'd 8992: out = 14'h1D27;
            14'd 8993: out = 14'h1D26;
            14'd 8994: out = 14'h1D26;
            14'd 8995: out = 14'h1D25;
            14'd 8996: out = 14'h1D24;
            14'd 8997: out = 14'h1D23;
            14'd 8998: out = 14'h1D22;
            14'd 8999: out = 14'h1D21;
            14'd 9000: out = 14'h1D21;
            14'd 9001: out = 14'h1D20;
            14'd 9002: out = 14'h1D1F;
            14'd 9003: out = 14'h1D1E;
            14'd 9004: out = 14'h1D1D;
            14'd 9005: out = 14'h1D1C;
            14'd 9006: out = 14'h1D1C;
            14'd 9007: out = 14'h1D1B;
            14'd 9008: out = 14'h1D1A;
            14'd 9009: out = 14'h1D19;
            14'd 9010: out = 14'h1D18;
            14'd 9011: out = 14'h1D17;
            14'd 9012: out = 14'h1D17;
            14'd 9013: out = 14'h1D16;
            14'd 9014: out = 14'h1D15;
            14'd 9015: out = 14'h1D14;
            14'd 9016: out = 14'h1D13;
            14'd 9017: out = 14'h1D12;
            14'd 9018: out = 14'h1D12;
            14'd 9019: out = 14'h1D11;
            14'd 9020: out = 14'h1D10;
            14'd 9021: out = 14'h1D0F;
            14'd 9022: out = 14'h1D0E;
            14'd 9023: out = 14'h1D0E;
            14'd 9024: out = 14'h1D0D;
            14'd 9025: out = 14'h1D0C;
            14'd 9026: out = 14'h1D0B;
            14'd 9027: out = 14'h1D0A;
            14'd 9028: out = 14'h1D09;
            14'd 9029: out = 14'h1D09;
            14'd 9030: out = 14'h1D08;
            14'd 9031: out = 14'h1D07;
            14'd 9032: out = 14'h1D06;
            14'd 9033: out = 14'h1D05;
            14'd 9034: out = 14'h1D04;
            14'd 9035: out = 14'h1D04;
            14'd 9036: out = 14'h1D03;
            14'd 9037: out = 14'h1D02;
            14'd 9038: out = 14'h1D01;
            14'd 9039: out = 14'h1D00;
            14'd 9040: out = 14'h1D00;
            14'd 9041: out = 14'h1CFF;
            14'd 9042: out = 14'h1CFE;
            14'd 9043: out = 14'h1CFD;
            14'd 9044: out = 14'h1CFC;
            14'd 9045: out = 14'h1CFB;
            14'd 9046: out = 14'h1CFB;
            14'd 9047: out = 14'h1CFA;
            14'd 9048: out = 14'h1CF9;
            14'd 9049: out = 14'h1CF8;
            14'd 9050: out = 14'h1CF7;
            14'd 9051: out = 14'h1CF7;
            14'd 9052: out = 14'h1CF6;
            14'd 9053: out = 14'h1CF5;
            14'd 9054: out = 14'h1CF4;
            14'd 9055: out = 14'h1CF3;
            14'd 9056: out = 14'h1CF2;
            14'd 9057: out = 14'h1CF2;
            14'd 9058: out = 14'h1CF1;
            14'd 9059: out = 14'h1CF0;
            14'd 9060: out = 14'h1CEF;
            14'd 9061: out = 14'h1CEE;
            14'd 9062: out = 14'h1CEE;
            14'd 9063: out = 14'h1CED;
            14'd 9064: out = 14'h1CEC;
            14'd 9065: out = 14'h1CEB;
            14'd 9066: out = 14'h1CEA;
            14'd 9067: out = 14'h1CE9;
            14'd 9068: out = 14'h1CE9;
            14'd 9069: out = 14'h1CE8;
            14'd 9070: out = 14'h1CE7;
            14'd 9071: out = 14'h1CE6;
            14'd 9072: out = 14'h1CE5;
            14'd 9073: out = 14'h1CE5;
            14'd 9074: out = 14'h1CE4;
            14'd 9075: out = 14'h1CE3;
            14'd 9076: out = 14'h1CE2;
            14'd 9077: out = 14'h1CE1;
            14'd 9078: out = 14'h1CE0;
            14'd 9079: out = 14'h1CE0;
            14'd 9080: out = 14'h1CDF;
            14'd 9081: out = 14'h1CDE;
            14'd 9082: out = 14'h1CDD;
            14'd 9083: out = 14'h1CDC;
            14'd 9084: out = 14'h1CDC;
            14'd 9085: out = 14'h1CDB;
            14'd 9086: out = 14'h1CDA;
            14'd 9087: out = 14'h1CD9;
            14'd 9088: out = 14'h1CD8;
            14'd 9089: out = 14'h1CD8;
            14'd 9090: out = 14'h1CD7;
            14'd 9091: out = 14'h1CD6;
            14'd 9092: out = 14'h1CD5;
            14'd 9093: out = 14'h1CD4;
            14'd 9094: out = 14'h1CD3;
            14'd 9095: out = 14'h1CD3;
            14'd 9096: out = 14'h1CD2;
            14'd 9097: out = 14'h1CD1;
            14'd 9098: out = 14'h1CD0;
            14'd 9099: out = 14'h1CCF;
            14'd 9100: out = 14'h1CCF;
            14'd 9101: out = 14'h1CCE;
            14'd 9102: out = 14'h1CCD;
            14'd 9103: out = 14'h1CCC;
            14'd 9104: out = 14'h1CCB;
            14'd 9105: out = 14'h1CCB;
            14'd 9106: out = 14'h1CCA;
            14'd 9107: out = 14'h1CC9;
            14'd 9108: out = 14'h1CC8;
            14'd 9109: out = 14'h1CC7;
            14'd 9110: out = 14'h1CC7;
            14'd 9111: out = 14'h1CC6;
            14'd 9112: out = 14'h1CC5;
            14'd 9113: out = 14'h1CC4;
            14'd 9114: out = 14'h1CC3;
            14'd 9115: out = 14'h1CC2;
            14'd 9116: out = 14'h1CC2;
            14'd 9117: out = 14'h1CC1;
            14'd 9118: out = 14'h1CC0;
            14'd 9119: out = 14'h1CBF;
            14'd 9120: out = 14'h1CBE;
            14'd 9121: out = 14'h1CBE;
            14'd 9122: out = 14'h1CBD;
            14'd 9123: out = 14'h1CBC;
            14'd 9124: out = 14'h1CBB;
            14'd 9125: out = 14'h1CBA;
            14'd 9126: out = 14'h1CBA;
            14'd 9127: out = 14'h1CB9;
            14'd 9128: out = 14'h1CB8;
            14'd 9129: out = 14'h1CB7;
            14'd 9130: out = 14'h1CB6;
            14'd 9131: out = 14'h1CB6;
            14'd 9132: out = 14'h1CB5;
            14'd 9133: out = 14'h1CB4;
            14'd 9134: out = 14'h1CB3;
            14'd 9135: out = 14'h1CB2;
            14'd 9136: out = 14'h1CB2;
            14'd 9137: out = 14'h1CB1;
            14'd 9138: out = 14'h1CB0;
            14'd 9139: out = 14'h1CAF;
            14'd 9140: out = 14'h1CAE;
            14'd 9141: out = 14'h1CAE;
            14'd 9142: out = 14'h1CAD;
            14'd 9143: out = 14'h1CAC;
            14'd 9144: out = 14'h1CAB;
            14'd 9145: out = 14'h1CAA;
            14'd 9146: out = 14'h1CAA;
            14'd 9147: out = 14'h1CA9;
            14'd 9148: out = 14'h1CA8;
            14'd 9149: out = 14'h1CA7;
            14'd 9150: out = 14'h1CA6;
            14'd 9151: out = 14'h1CA6;
            14'd 9152: out = 14'h1CA5;
            14'd 9153: out = 14'h1CA4;
            14'd 9154: out = 14'h1CA3;
            14'd 9155: out = 14'h1CA2;
            14'd 9156: out = 14'h1CA1;
            14'd 9157: out = 14'h1CA1;
            14'd 9158: out = 14'h1CA0;
            14'd 9159: out = 14'h1C9F;
            14'd 9160: out = 14'h1C9E;
            14'd 9161: out = 14'h1C9D;
            14'd 9162: out = 14'h1C9D;
            14'd 9163: out = 14'h1C9C;
            14'd 9164: out = 14'h1C9B;
            14'd 9165: out = 14'h1C9A;
            14'd 9166: out = 14'h1C99;
            14'd 9167: out = 14'h1C99;
            14'd 9168: out = 14'h1C98;
            14'd 9169: out = 14'h1C97;
            14'd 9170: out = 14'h1C96;
            14'd 9171: out = 14'h1C96;
            14'd 9172: out = 14'h1C95;
            14'd 9173: out = 14'h1C94;
            14'd 9174: out = 14'h1C93;
            14'd 9175: out = 14'h1C92;
            14'd 9176: out = 14'h1C92;
            14'd 9177: out = 14'h1C91;
            14'd 9178: out = 14'h1C90;
            14'd 9179: out = 14'h1C8F;
            14'd 9180: out = 14'h1C8E;
            14'd 9181: out = 14'h1C8E;
            14'd 9182: out = 14'h1C8D;
            14'd 9183: out = 14'h1C8C;
            14'd 9184: out = 14'h1C8B;
            14'd 9185: out = 14'h1C8A;
            14'd 9186: out = 14'h1C8A;
            14'd 9187: out = 14'h1C89;
            14'd 9188: out = 14'h1C88;
            14'd 9189: out = 14'h1C87;
            14'd 9190: out = 14'h1C86;
            14'd 9191: out = 14'h1C86;
            14'd 9192: out = 14'h1C85;
            14'd 9193: out = 14'h1C84;
            14'd 9194: out = 14'h1C83;
            14'd 9195: out = 14'h1C82;
            14'd 9196: out = 14'h1C82;
            14'd 9197: out = 14'h1C81;
            14'd 9198: out = 14'h1C80;
            14'd 9199: out = 14'h1C7F;
            14'd 9200: out = 14'h1C7E;
            14'd 9201: out = 14'h1C7E;
            14'd 9202: out = 14'h1C7D;
            14'd 9203: out = 14'h1C7C;
            14'd 9204: out = 14'h1C7B;
            14'd 9205: out = 14'h1C7A;
            14'd 9206: out = 14'h1C7A;
            14'd 9207: out = 14'h1C79;
            14'd 9208: out = 14'h1C78;
            14'd 9209: out = 14'h1C77;
            14'd 9210: out = 14'h1C77;
            14'd 9211: out = 14'h1C76;
            14'd 9212: out = 14'h1C75;
            14'd 9213: out = 14'h1C74;
            14'd 9214: out = 14'h1C73;
            14'd 9215: out = 14'h1C73;
            14'd 9216: out = 14'h1C72;
            14'd 9217: out = 14'h1C71;
            14'd 9218: out = 14'h1C70;
            14'd 9219: out = 14'h1C6F;
            14'd 9220: out = 14'h1C6F;
            14'd 9221: out = 14'h1C6E;
            14'd 9222: out = 14'h1C6D;
            14'd 9223: out = 14'h1C6C;
            14'd 9224: out = 14'h1C6B;
            14'd 9225: out = 14'h1C6B;
            14'd 9226: out = 14'h1C6A;
            14'd 9227: out = 14'h1C69;
            14'd 9228: out = 14'h1C68;
            14'd 9229: out = 14'h1C68;
            14'd 9230: out = 14'h1C67;
            14'd 9231: out = 14'h1C66;
            14'd 9232: out = 14'h1C65;
            14'd 9233: out = 14'h1C64;
            14'd 9234: out = 14'h1C64;
            14'd 9235: out = 14'h1C63;
            14'd 9236: out = 14'h1C62;
            14'd 9237: out = 14'h1C61;
            14'd 9238: out = 14'h1C60;
            14'd 9239: out = 14'h1C60;
            14'd 9240: out = 14'h1C5F;
            14'd 9241: out = 14'h1C5E;
            14'd 9242: out = 14'h1C5D;
            14'd 9243: out = 14'h1C5D;
            14'd 9244: out = 14'h1C5C;
            14'd 9245: out = 14'h1C5B;
            14'd 9246: out = 14'h1C5A;
            14'd 9247: out = 14'h1C59;
            14'd 9248: out = 14'h1C59;
            14'd 9249: out = 14'h1C58;
            14'd 9250: out = 14'h1C57;
            14'd 9251: out = 14'h1C56;
            14'd 9252: out = 14'h1C55;
            14'd 9253: out = 14'h1C55;
            14'd 9254: out = 14'h1C54;
            14'd 9255: out = 14'h1C53;
            14'd 9256: out = 14'h1C52;
            14'd 9257: out = 14'h1C52;
            14'd 9258: out = 14'h1C51;
            14'd 9259: out = 14'h1C50;
            14'd 9260: out = 14'h1C4F;
            14'd 9261: out = 14'h1C4E;
            14'd 9262: out = 14'h1C4E;
            14'd 9263: out = 14'h1C4D;
            14'd 9264: out = 14'h1C4C;
            14'd 9265: out = 14'h1C4B;
            14'd 9266: out = 14'h1C4A;
            14'd 9267: out = 14'h1C4A;
            14'd 9268: out = 14'h1C49;
            14'd 9269: out = 14'h1C48;
            14'd 9270: out = 14'h1C47;
            14'd 9271: out = 14'h1C47;
            14'd 9272: out = 14'h1C46;
            14'd 9273: out = 14'h1C45;
            14'd 9274: out = 14'h1C44;
            14'd 9275: out = 14'h1C43;
            14'd 9276: out = 14'h1C43;
            14'd 9277: out = 14'h1C42;
            14'd 9278: out = 14'h1C41;
            14'd 9279: out = 14'h1C40;
            14'd 9280: out = 14'h1C40;
            14'd 9281: out = 14'h1C3F;
            14'd 9282: out = 14'h1C3E;
            14'd 9283: out = 14'h1C3D;
            14'd 9284: out = 14'h1C3C;
            14'd 9285: out = 14'h1C3C;
            14'd 9286: out = 14'h1C3B;
            14'd 9287: out = 14'h1C3A;
            14'd 9288: out = 14'h1C39;
            14'd 9289: out = 14'h1C39;
            14'd 9290: out = 14'h1C38;
            14'd 9291: out = 14'h1C37;
            14'd 9292: out = 14'h1C36;
            14'd 9293: out = 14'h1C35;
            14'd 9294: out = 14'h1C35;
            14'd 9295: out = 14'h1C34;
            14'd 9296: out = 14'h1C33;
            14'd 9297: out = 14'h1C32;
            14'd 9298: out = 14'h1C32;
            14'd 9299: out = 14'h1C31;
            14'd 9300: out = 14'h1C30;
            14'd 9301: out = 14'h1C2F;
            14'd 9302: out = 14'h1C2E;
            14'd 9303: out = 14'h1C2E;
            14'd 9304: out = 14'h1C2D;
            14'd 9305: out = 14'h1C2C;
            14'd 9306: out = 14'h1C2B;
            14'd 9307: out = 14'h1C2B;
            14'd 9308: out = 14'h1C2A;
            14'd 9309: out = 14'h1C29;
            14'd 9310: out = 14'h1C28;
            14'd 9311: out = 14'h1C27;
            14'd 9312: out = 14'h1C27;
            14'd 9313: out = 14'h1C26;
            14'd 9314: out = 14'h1C25;
            14'd 9315: out = 14'h1C24;
            14'd 9316: out = 14'h1C24;
            14'd 9317: out = 14'h1C23;
            14'd 9318: out = 14'h1C22;
            14'd 9319: out = 14'h1C21;
            14'd 9320: out = 14'h1C21;
            14'd 9321: out = 14'h1C20;
            14'd 9322: out = 14'h1C1F;
            14'd 9323: out = 14'h1C1E;
            14'd 9324: out = 14'h1C1D;
            14'd 9325: out = 14'h1C1D;
            14'd 9326: out = 14'h1C1C;
            14'd 9327: out = 14'h1C1B;
            14'd 9328: out = 14'h1C1A;
            14'd 9329: out = 14'h1C1A;
            14'd 9330: out = 14'h1C19;
            14'd 9331: out = 14'h1C18;
            14'd 9332: out = 14'h1C17;
            14'd 9333: out = 14'h1C16;
            14'd 9334: out = 14'h1C16;
            14'd 9335: out = 14'h1C15;
            14'd 9336: out = 14'h1C14;
            14'd 9337: out = 14'h1C13;
            14'd 9338: out = 14'h1C13;
            14'd 9339: out = 14'h1C12;
            14'd 9340: out = 14'h1C11;
            14'd 9341: out = 14'h1C10;
            14'd 9342: out = 14'h1C10;
            14'd 9343: out = 14'h1C0F;
            14'd 9344: out = 14'h1C0E;
            14'd 9345: out = 14'h1C0D;
            14'd 9346: out = 14'h1C0C;
            14'd 9347: out = 14'h1C0C;
            14'd 9348: out = 14'h1C0B;
            14'd 9349: out = 14'h1C0A;
            14'd 9350: out = 14'h1C09;
            14'd 9351: out = 14'h1C09;
            14'd 9352: out = 14'h1C08;
            14'd 9353: out = 14'h1C07;
            14'd 9354: out = 14'h1C06;
            14'd 9355: out = 14'h1C06;
            14'd 9356: out = 14'h1C05;
            14'd 9357: out = 14'h1C04;
            14'd 9358: out = 14'h1C03;
            14'd 9359: out = 14'h1C03;
            14'd 9360: out = 14'h1C02;
            14'd 9361: out = 14'h1C01;
            14'd 9362: out = 14'h1C00;
            14'd 9363: out = 14'h1BFF;
            14'd 9364: out = 14'h1BFF;
            14'd 9365: out = 14'h1BFE;
            14'd 9366: out = 14'h1BFD;
            14'd 9367: out = 14'h1BFC;
            14'd 9368: out = 14'h1BFC;
            14'd 9369: out = 14'h1BFB;
            14'd 9370: out = 14'h1BFA;
            14'd 9371: out = 14'h1BF9;
            14'd 9372: out = 14'h1BF9;
            14'd 9373: out = 14'h1BF8;
            14'd 9374: out = 14'h1BF7;
            14'd 9375: out = 14'h1BF6;
            14'd 9376: out = 14'h1BF6;
            14'd 9377: out = 14'h1BF5;
            14'd 9378: out = 14'h1BF4;
            14'd 9379: out = 14'h1BF3;
            14'd 9380: out = 14'h1BF2;
            14'd 9381: out = 14'h1BF2;
            14'd 9382: out = 14'h1BF1;
            14'd 9383: out = 14'h1BF0;
            14'd 9384: out = 14'h1BEF;
            14'd 9385: out = 14'h1BEF;
            14'd 9386: out = 14'h1BEE;
            14'd 9387: out = 14'h1BED;
            14'd 9388: out = 14'h1BEC;
            14'd 9389: out = 14'h1BEC;
            14'd 9390: out = 14'h1BEB;
            14'd 9391: out = 14'h1BEA;
            14'd 9392: out = 14'h1BE9;
            14'd 9393: out = 14'h1BE9;
            14'd 9394: out = 14'h1BE8;
            14'd 9395: out = 14'h1BE7;
            14'd 9396: out = 14'h1BE6;
            14'd 9397: out = 14'h1BE6;
            14'd 9398: out = 14'h1BE5;
            14'd 9399: out = 14'h1BE4;
            14'd 9400: out = 14'h1BE3;
            14'd 9401: out = 14'h1BE2;
            14'd 9402: out = 14'h1BE2;
            14'd 9403: out = 14'h1BE1;
            14'd 9404: out = 14'h1BE0;
            14'd 9405: out = 14'h1BDF;
            14'd 9406: out = 14'h1BDF;
            14'd 9407: out = 14'h1BDE;
            14'd 9408: out = 14'h1BDD;
            14'd 9409: out = 14'h1BDC;
            14'd 9410: out = 14'h1BDC;
            14'd 9411: out = 14'h1BDB;
            14'd 9412: out = 14'h1BDA;
            14'd 9413: out = 14'h1BD9;
            14'd 9414: out = 14'h1BD9;
            14'd 9415: out = 14'h1BD8;
            14'd 9416: out = 14'h1BD7;
            14'd 9417: out = 14'h1BD6;
            14'd 9418: out = 14'h1BD6;
            14'd 9419: out = 14'h1BD5;
            14'd 9420: out = 14'h1BD4;
            14'd 9421: out = 14'h1BD3;
            14'd 9422: out = 14'h1BD3;
            14'd 9423: out = 14'h1BD2;
            14'd 9424: out = 14'h1BD1;
            14'd 9425: out = 14'h1BD0;
            14'd 9426: out = 14'h1BD0;
            14'd 9427: out = 14'h1BCF;
            14'd 9428: out = 14'h1BCE;
            14'd 9429: out = 14'h1BCD;
            14'd 9430: out = 14'h1BCD;
            14'd 9431: out = 14'h1BCC;
            14'd 9432: out = 14'h1BCB;
            14'd 9433: out = 14'h1BCA;
            14'd 9434: out = 14'h1BCA;
            14'd 9435: out = 14'h1BC9;
            14'd 9436: out = 14'h1BC8;
            14'd 9437: out = 14'h1BC7;
            14'd 9438: out = 14'h1BC6;
            14'd 9439: out = 14'h1BC6;
            14'd 9440: out = 14'h1BC5;
            14'd 9441: out = 14'h1BC4;
            14'd 9442: out = 14'h1BC3;
            14'd 9443: out = 14'h1BC3;
            14'd 9444: out = 14'h1BC2;
            14'd 9445: out = 14'h1BC1;
            14'd 9446: out = 14'h1BC0;
            14'd 9447: out = 14'h1BC0;
            14'd 9448: out = 14'h1BBF;
            14'd 9449: out = 14'h1BBE;
            14'd 9450: out = 14'h1BBD;
            14'd 9451: out = 14'h1BBD;
            14'd 9452: out = 14'h1BBC;
            14'd 9453: out = 14'h1BBB;
            14'd 9454: out = 14'h1BBA;
            14'd 9455: out = 14'h1BBA;
            14'd 9456: out = 14'h1BB9;
            14'd 9457: out = 14'h1BB8;
            14'd 9458: out = 14'h1BB7;
            14'd 9459: out = 14'h1BB7;
            14'd 9460: out = 14'h1BB6;
            14'd 9461: out = 14'h1BB5;
            14'd 9462: out = 14'h1BB4;
            14'd 9463: out = 14'h1BB4;
            14'd 9464: out = 14'h1BB3;
            14'd 9465: out = 14'h1BB2;
            14'd 9466: out = 14'h1BB1;
            14'd 9467: out = 14'h1BB1;
            14'd 9468: out = 14'h1BB0;
            14'd 9469: out = 14'h1BAF;
            14'd 9470: out = 14'h1BAE;
            14'd 9471: out = 14'h1BAE;
            14'd 9472: out = 14'h1BAD;
            14'd 9473: out = 14'h1BAC;
            14'd 9474: out = 14'h1BAB;
            14'd 9475: out = 14'h1BAB;
            14'd 9476: out = 14'h1BAA;
            14'd 9477: out = 14'h1BA9;
            14'd 9478: out = 14'h1BA8;
            14'd 9479: out = 14'h1BA8;
            14'd 9480: out = 14'h1BA7;
            14'd 9481: out = 14'h1BA6;
            14'd 9482: out = 14'h1BA6;
            14'd 9483: out = 14'h1BA5;
            14'd 9484: out = 14'h1BA4;
            14'd 9485: out = 14'h1BA3;
            14'd 9486: out = 14'h1BA3;
            14'd 9487: out = 14'h1BA2;
            14'd 9488: out = 14'h1BA1;
            14'd 9489: out = 14'h1BA0;
            14'd 9490: out = 14'h1BA0;
            14'd 9491: out = 14'h1B9F;
            14'd 9492: out = 14'h1B9E;
            14'd 9493: out = 14'h1B9D;
            14'd 9494: out = 14'h1B9D;
            14'd 9495: out = 14'h1B9C;
            14'd 9496: out = 14'h1B9B;
            14'd 9497: out = 14'h1B9A;
            14'd 9498: out = 14'h1B9A;
            14'd 9499: out = 14'h1B99;
            14'd 9500: out = 14'h1B98;
            14'd 9501: out = 14'h1B97;
            14'd 9502: out = 14'h1B97;
            14'd 9503: out = 14'h1B96;
            14'd 9504: out = 14'h1B95;
            14'd 9505: out = 14'h1B94;
            14'd 9506: out = 14'h1B94;
            14'd 9507: out = 14'h1B93;
            14'd 9508: out = 14'h1B92;
            14'd 9509: out = 14'h1B91;
            14'd 9510: out = 14'h1B91;
            14'd 9511: out = 14'h1B90;
            14'd 9512: out = 14'h1B8F;
            14'd 9513: out = 14'h1B8E;
            14'd 9514: out = 14'h1B8E;
            14'd 9515: out = 14'h1B8D;
            14'd 9516: out = 14'h1B8C;
            14'd 9517: out = 14'h1B8B;
            14'd 9518: out = 14'h1B8B;
            14'd 9519: out = 14'h1B8A;
            14'd 9520: out = 14'h1B89;
            14'd 9521: out = 14'h1B89;
            14'd 9522: out = 14'h1B88;
            14'd 9523: out = 14'h1B87;
            14'd 9524: out = 14'h1B86;
            14'd 9525: out = 14'h1B86;
            14'd 9526: out = 14'h1B85;
            14'd 9527: out = 14'h1B84;
            14'd 9528: out = 14'h1B83;
            14'd 9529: out = 14'h1B83;
            14'd 9530: out = 14'h1B82;
            14'd 9531: out = 14'h1B81;
            14'd 9532: out = 14'h1B80;
            14'd 9533: out = 14'h1B80;
            14'd 9534: out = 14'h1B7F;
            14'd 9535: out = 14'h1B7E;
            14'd 9536: out = 14'h1B7D;
            14'd 9537: out = 14'h1B7D;
            14'd 9538: out = 14'h1B7C;
            14'd 9539: out = 14'h1B7B;
            14'd 9540: out = 14'h1B7A;
            14'd 9541: out = 14'h1B7A;
            14'd 9542: out = 14'h1B79;
            14'd 9543: out = 14'h1B78;
            14'd 9544: out = 14'h1B78;
            14'd 9545: out = 14'h1B77;
            14'd 9546: out = 14'h1B76;
            14'd 9547: out = 14'h1B75;
            14'd 9548: out = 14'h1B75;
            14'd 9549: out = 14'h1B74;
            14'd 9550: out = 14'h1B73;
            14'd 9551: out = 14'h1B72;
            14'd 9552: out = 14'h1B72;
            14'd 9553: out = 14'h1B71;
            14'd 9554: out = 14'h1B70;
            14'd 9555: out = 14'h1B6F;
            14'd 9556: out = 14'h1B6F;
            14'd 9557: out = 14'h1B6E;
            14'd 9558: out = 14'h1B6D;
            14'd 9559: out = 14'h1B6C;
            14'd 9560: out = 14'h1B6C;
            14'd 9561: out = 14'h1B6B;
            14'd 9562: out = 14'h1B6A;
            14'd 9563: out = 14'h1B6A;
            14'd 9564: out = 14'h1B69;
            14'd 9565: out = 14'h1B68;
            14'd 9566: out = 14'h1B67;
            14'd 9567: out = 14'h1B67;
            14'd 9568: out = 14'h1B66;
            14'd 9569: out = 14'h1B65;
            14'd 9570: out = 14'h1B64;
            14'd 9571: out = 14'h1B64;
            14'd 9572: out = 14'h1B63;
            14'd 9573: out = 14'h1B62;
            14'd 9574: out = 14'h1B61;
            14'd 9575: out = 14'h1B61;
            14'd 9576: out = 14'h1B60;
            14'd 9577: out = 14'h1B5F;
            14'd 9578: out = 14'h1B5F;
            14'd 9579: out = 14'h1B5E;
            14'd 9580: out = 14'h1B5D;
            14'd 9581: out = 14'h1B5C;
            14'd 9582: out = 14'h1B5C;
            14'd 9583: out = 14'h1B5B;
            14'd 9584: out = 14'h1B5A;
            14'd 9585: out = 14'h1B59;
            14'd 9586: out = 14'h1B59;
            14'd 9587: out = 14'h1B58;
            14'd 9588: out = 14'h1B57;
            14'd 9589: out = 14'h1B57;
            14'd 9590: out = 14'h1B56;
            14'd 9591: out = 14'h1B55;
            14'd 9592: out = 14'h1B54;
            14'd 9593: out = 14'h1B54;
            14'd 9594: out = 14'h1B53;
            14'd 9595: out = 14'h1B52;
            14'd 9596: out = 14'h1B51;
            14'd 9597: out = 14'h1B51;
            14'd 9598: out = 14'h1B50;
            14'd 9599: out = 14'h1B4F;
            14'd 9600: out = 14'h1B4F;
            14'd 9601: out = 14'h1B4E;
            14'd 9602: out = 14'h1B4D;
            14'd 9603: out = 14'h1B4C;
            14'd 9604: out = 14'h1B4C;
            14'd 9605: out = 14'h1B4B;
            14'd 9606: out = 14'h1B4A;
            14'd 9607: out = 14'h1B49;
            14'd 9608: out = 14'h1B49;
            14'd 9609: out = 14'h1B48;
            14'd 9610: out = 14'h1B47;
            14'd 9611: out = 14'h1B47;
            14'd 9612: out = 14'h1B46;
            14'd 9613: out = 14'h1B45;
            14'd 9614: out = 14'h1B44;
            14'd 9615: out = 14'h1B44;
            14'd 9616: out = 14'h1B43;
            14'd 9617: out = 14'h1B42;
            14'd 9618: out = 14'h1B41;
            14'd 9619: out = 14'h1B41;
            14'd 9620: out = 14'h1B40;
            14'd 9621: out = 14'h1B3F;
            14'd 9622: out = 14'h1B3F;
            14'd 9623: out = 14'h1B3E;
            14'd 9624: out = 14'h1B3D;
            14'd 9625: out = 14'h1B3C;
            14'd 9626: out = 14'h1B3C;
            14'd 9627: out = 14'h1B3B;
            14'd 9628: out = 14'h1B3A;
            14'd 9629: out = 14'h1B39;
            14'd 9630: out = 14'h1B39;
            14'd 9631: out = 14'h1B38;
            14'd 9632: out = 14'h1B37;
            14'd 9633: out = 14'h1B37;
            14'd 9634: out = 14'h1B36;
            14'd 9635: out = 14'h1B35;
            14'd 9636: out = 14'h1B34;
            14'd 9637: out = 14'h1B34;
            14'd 9638: out = 14'h1B33;
            14'd 9639: out = 14'h1B32;
            14'd 9640: out = 14'h1B32;
            14'd 9641: out = 14'h1B31;
            14'd 9642: out = 14'h1B30;
            14'd 9643: out = 14'h1B2F;
            14'd 9644: out = 14'h1B2F;
            14'd 9645: out = 14'h1B2E;
            14'd 9646: out = 14'h1B2D;
            14'd 9647: out = 14'h1B2C;
            14'd 9648: out = 14'h1B2C;
            14'd 9649: out = 14'h1B2B;
            14'd 9650: out = 14'h1B2A;
            14'd 9651: out = 14'h1B2A;
            14'd 9652: out = 14'h1B29;
            14'd 9653: out = 14'h1B28;
            14'd 9654: out = 14'h1B27;
            14'd 9655: out = 14'h1B27;
            14'd 9656: out = 14'h1B26;
            14'd 9657: out = 14'h1B25;
            14'd 9658: out = 14'h1B25;
            14'd 9659: out = 14'h1B24;
            14'd 9660: out = 14'h1B23;
            14'd 9661: out = 14'h1B22;
            14'd 9662: out = 14'h1B22;
            14'd 9663: out = 14'h1B21;
            14'd 9664: out = 14'h1B20;
            14'd 9665: out = 14'h1B1F;
            14'd 9666: out = 14'h1B1F;
            14'd 9667: out = 14'h1B1E;
            14'd 9668: out = 14'h1B1D;
            14'd 9669: out = 14'h1B1D;
            14'd 9670: out = 14'h1B1C;
            14'd 9671: out = 14'h1B1B;
            14'd 9672: out = 14'h1B1A;
            14'd 9673: out = 14'h1B1A;
            14'd 9674: out = 14'h1B19;
            14'd 9675: out = 14'h1B18;
            14'd 9676: out = 14'h1B18;
            14'd 9677: out = 14'h1B17;
            14'd 9678: out = 14'h1B16;
            14'd 9679: out = 14'h1B15;
            14'd 9680: out = 14'h1B15;
            14'd 9681: out = 14'h1B14;
            14'd 9682: out = 14'h1B13;
            14'd 9683: out = 14'h1B13;
            14'd 9684: out = 14'h1B12;
            14'd 9685: out = 14'h1B11;
            14'd 9686: out = 14'h1B10;
            14'd 9687: out = 14'h1B10;
            14'd 9688: out = 14'h1B0F;
            14'd 9689: out = 14'h1B0E;
            14'd 9690: out = 14'h1B0E;
            14'd 9691: out = 14'h1B0D;
            14'd 9692: out = 14'h1B0C;
            14'd 9693: out = 14'h1B0B;
            14'd 9694: out = 14'h1B0B;
            14'd 9695: out = 14'h1B0A;
            14'd 9696: out = 14'h1B09;
            14'd 9697: out = 14'h1B09;
            14'd 9698: out = 14'h1B08;
            14'd 9699: out = 14'h1B07;
            14'd 9700: out = 14'h1B06;
            14'd 9701: out = 14'h1B06;
            14'd 9702: out = 14'h1B05;
            14'd 9703: out = 14'h1B04;
            14'd 9704: out = 14'h1B04;
            14'd 9705: out = 14'h1B03;
            14'd 9706: out = 14'h1B02;
            14'd 9707: out = 14'h1B01;
            14'd 9708: out = 14'h1B01;
            14'd 9709: out = 14'h1B00;
            14'd 9710: out = 14'h1AFF;
            14'd 9711: out = 14'h1AFF;
            14'd 9712: out = 14'h1AFE;
            14'd 9713: out = 14'h1AFD;
            14'd 9714: out = 14'h1AFC;
            14'd 9715: out = 14'h1AFC;
            14'd 9716: out = 14'h1AFB;
            14'd 9717: out = 14'h1AFA;
            14'd 9718: out = 14'h1AFA;
            14'd 9719: out = 14'h1AF9;
            14'd 9720: out = 14'h1AF8;
            14'd 9721: out = 14'h1AF7;
            14'd 9722: out = 14'h1AF7;
            14'd 9723: out = 14'h1AF6;
            14'd 9724: out = 14'h1AF5;
            14'd 9725: out = 14'h1AF5;
            14'd 9726: out = 14'h1AF4;
            14'd 9727: out = 14'h1AF3;
            14'd 9728: out = 14'h1AF3;
            14'd 9729: out = 14'h1AF2;
            14'd 9730: out = 14'h1AF1;
            14'd 9731: out = 14'h1AF0;
            14'd 9732: out = 14'h1AF0;
            14'd 9733: out = 14'h1AEF;
            14'd 9734: out = 14'h1AEE;
            14'd 9735: out = 14'h1AEE;
            14'd 9736: out = 14'h1AED;
            14'd 9737: out = 14'h1AEC;
            14'd 9738: out = 14'h1AEB;
            14'd 9739: out = 14'h1AEB;
            14'd 9740: out = 14'h1AEA;
            14'd 9741: out = 14'h1AE9;
            14'd 9742: out = 14'h1AE9;
            14'd 9743: out = 14'h1AE8;
            14'd 9744: out = 14'h1AE7;
            14'd 9745: out = 14'h1AE6;
            14'd 9746: out = 14'h1AE6;
            14'd 9747: out = 14'h1AE5;
            14'd 9748: out = 14'h1AE4;
            14'd 9749: out = 14'h1AE4;
            14'd 9750: out = 14'h1AE3;
            14'd 9751: out = 14'h1AE2;
            14'd 9752: out = 14'h1AE2;
            14'd 9753: out = 14'h1AE1;
            14'd 9754: out = 14'h1AE0;
            14'd 9755: out = 14'h1ADF;
            14'd 9756: out = 14'h1ADF;
            14'd 9757: out = 14'h1ADE;
            14'd 9758: out = 14'h1ADD;
            14'd 9759: out = 14'h1ADD;
            14'd 9760: out = 14'h1ADC;
            14'd 9761: out = 14'h1ADB;
            14'd 9762: out = 14'h1ADA;
            14'd 9763: out = 14'h1ADA;
            14'd 9764: out = 14'h1AD9;
            14'd 9765: out = 14'h1AD8;
            14'd 9766: out = 14'h1AD8;
            14'd 9767: out = 14'h1AD7;
            14'd 9768: out = 14'h1AD6;
            14'd 9769: out = 14'h1AD6;
            14'd 9770: out = 14'h1AD5;
            14'd 9771: out = 14'h1AD4;
            14'd 9772: out = 14'h1AD3;
            14'd 9773: out = 14'h1AD3;
            14'd 9774: out = 14'h1AD2;
            14'd 9775: out = 14'h1AD1;
            14'd 9776: out = 14'h1AD1;
            14'd 9777: out = 14'h1AD0;
            14'd 9778: out = 14'h1ACF;
            14'd 9779: out = 14'h1ACF;
            14'd 9780: out = 14'h1ACE;
            14'd 9781: out = 14'h1ACD;
            14'd 9782: out = 14'h1ACC;
            14'd 9783: out = 14'h1ACC;
            14'd 9784: out = 14'h1ACB;
            14'd 9785: out = 14'h1ACA;
            14'd 9786: out = 14'h1ACA;
            14'd 9787: out = 14'h1AC9;
            14'd 9788: out = 14'h1AC8;
            14'd 9789: out = 14'h1AC8;
            14'd 9790: out = 14'h1AC7;
            14'd 9791: out = 14'h1AC6;
            14'd 9792: out = 14'h1AC5;
            14'd 9793: out = 14'h1AC5;
            14'd 9794: out = 14'h1AC4;
            14'd 9795: out = 14'h1AC3;
            14'd 9796: out = 14'h1AC3;
            14'd 9797: out = 14'h1AC2;
            14'd 9798: out = 14'h1AC1;
            14'd 9799: out = 14'h1AC1;
            14'd 9800: out = 14'h1AC0;
            14'd 9801: out = 14'h1ABF;
            14'd 9802: out = 14'h1ABE;
            14'd 9803: out = 14'h1ABE;
            14'd 9804: out = 14'h1ABD;
            14'd 9805: out = 14'h1ABC;
            14'd 9806: out = 14'h1ABC;
            14'd 9807: out = 14'h1ABB;
            14'd 9808: out = 14'h1ABA;
            14'd 9809: out = 14'h1ABA;
            14'd 9810: out = 14'h1AB9;
            14'd 9811: out = 14'h1AB8;
            14'd 9812: out = 14'h1AB7;
            14'd 9813: out = 14'h1AB7;
            14'd 9814: out = 14'h1AB6;
            14'd 9815: out = 14'h1AB5;
            14'd 9816: out = 14'h1AB5;
            14'd 9817: out = 14'h1AB4;
            14'd 9818: out = 14'h1AB3;
            14'd 9819: out = 14'h1AB3;
            14'd 9820: out = 14'h1AB2;
            14'd 9821: out = 14'h1AB1;
            14'd 9822: out = 14'h1AB1;
            14'd 9823: out = 14'h1AB0;
            14'd 9824: out = 14'h1AAF;
            14'd 9825: out = 14'h1AAE;
            14'd 9826: out = 14'h1AAE;
            14'd 9827: out = 14'h1AAD;
            14'd 9828: out = 14'h1AAC;
            14'd 9829: out = 14'h1AAC;
            14'd 9830: out = 14'h1AAB;
            14'd 9831: out = 14'h1AAA;
            14'd 9832: out = 14'h1AAA;
            14'd 9833: out = 14'h1AA9;
            14'd 9834: out = 14'h1AA8;
            14'd 9835: out = 14'h1AA7;
            14'd 9836: out = 14'h1AA7;
            14'd 9837: out = 14'h1AA6;
            14'd 9838: out = 14'h1AA5;
            14'd 9839: out = 14'h1AA5;
            14'd 9840: out = 14'h1AA4;
            14'd 9841: out = 14'h1AA3;
            14'd 9842: out = 14'h1AA3;
            14'd 9843: out = 14'h1AA2;
            14'd 9844: out = 14'h1AA1;
            14'd 9845: out = 14'h1AA1;
            14'd 9846: out = 14'h1AA0;
            14'd 9847: out = 14'h1A9F;
            14'd 9848: out = 14'h1A9E;
            14'd 9849: out = 14'h1A9E;
            14'd 9850: out = 14'h1A9D;
            14'd 9851: out = 14'h1A9C;
            14'd 9852: out = 14'h1A9C;
            14'd 9853: out = 14'h1A9B;
            14'd 9854: out = 14'h1A9A;
            14'd 9855: out = 14'h1A9A;
            14'd 9856: out = 14'h1A99;
            14'd 9857: out = 14'h1A98;
            14'd 9858: out = 14'h1A98;
            14'd 9859: out = 14'h1A97;
            14'd 9860: out = 14'h1A96;
            14'd 9861: out = 14'h1A95;
            14'd 9862: out = 14'h1A95;
            14'd 9863: out = 14'h1A94;
            14'd 9864: out = 14'h1A93;
            14'd 9865: out = 14'h1A93;
            14'd 9866: out = 14'h1A92;
            14'd 9867: out = 14'h1A91;
            14'd 9868: out = 14'h1A91;
            14'd 9869: out = 14'h1A90;
            14'd 9870: out = 14'h1A8F;
            14'd 9871: out = 14'h1A8F;
            14'd 9872: out = 14'h1A8E;
            14'd 9873: out = 14'h1A8D;
            14'd 9874: out = 14'h1A8D;
            14'd 9875: out = 14'h1A8C;
            14'd 9876: out = 14'h1A8B;
            14'd 9877: out = 14'h1A8A;
            14'd 9878: out = 14'h1A8A;
            14'd 9879: out = 14'h1A89;
            14'd 9880: out = 14'h1A88;
            14'd 9881: out = 14'h1A88;
            14'd 9882: out = 14'h1A87;
            14'd 9883: out = 14'h1A86;
            14'd 9884: out = 14'h1A86;
            14'd 9885: out = 14'h1A85;
            14'd 9886: out = 14'h1A84;
            14'd 9887: out = 14'h1A84;
            14'd 9888: out = 14'h1A83;
            14'd 9889: out = 14'h1A82;
            14'd 9890: out = 14'h1A82;
            14'd 9891: out = 14'h1A81;
            14'd 9892: out = 14'h1A80;
            14'd 9893: out = 14'h1A7F;
            14'd 9894: out = 14'h1A7F;
            14'd 9895: out = 14'h1A7E;
            14'd 9896: out = 14'h1A7D;
            14'd 9897: out = 14'h1A7D;
            14'd 9898: out = 14'h1A7C;
            14'd 9899: out = 14'h1A7B;
            14'd 9900: out = 14'h1A7B;
            14'd 9901: out = 14'h1A7A;
            14'd 9902: out = 14'h1A79;
            14'd 9903: out = 14'h1A79;
            14'd 9904: out = 14'h1A78;
            14'd 9905: out = 14'h1A77;
            14'd 9906: out = 14'h1A77;
            14'd 9907: out = 14'h1A76;
            14'd 9908: out = 14'h1A75;
            14'd 9909: out = 14'h1A75;
            14'd 9910: out = 14'h1A74;
            14'd 9911: out = 14'h1A73;
            14'd 9912: out = 14'h1A72;
            14'd 9913: out = 14'h1A72;
            14'd 9914: out = 14'h1A71;
            14'd 9915: out = 14'h1A70;
            14'd 9916: out = 14'h1A70;
            14'd 9917: out = 14'h1A6F;
            14'd 9918: out = 14'h1A6E;
            14'd 9919: out = 14'h1A6E;
            14'd 9920: out = 14'h1A6D;
            14'd 9921: out = 14'h1A6C;
            14'd 9922: out = 14'h1A6C;
            14'd 9923: out = 14'h1A6B;
            14'd 9924: out = 14'h1A6A;
            14'd 9925: out = 14'h1A6A;
            14'd 9926: out = 14'h1A69;
            14'd 9927: out = 14'h1A68;
            14'd 9928: out = 14'h1A68;
            14'd 9929: out = 14'h1A67;
            14'd 9930: out = 14'h1A66;
            14'd 9931: out = 14'h1A66;
            14'd 9932: out = 14'h1A65;
            14'd 9933: out = 14'h1A64;
            14'd 9934: out = 14'h1A63;
            14'd 9935: out = 14'h1A63;
            14'd 9936: out = 14'h1A62;
            14'd 9937: out = 14'h1A61;
            14'd 9938: out = 14'h1A61;
            14'd 9939: out = 14'h1A60;
            14'd 9940: out = 14'h1A5F;
            14'd 9941: out = 14'h1A5F;
            14'd 9942: out = 14'h1A5E;
            14'd 9943: out = 14'h1A5D;
            14'd 9944: out = 14'h1A5D;
            14'd 9945: out = 14'h1A5C;
            14'd 9946: out = 14'h1A5B;
            14'd 9947: out = 14'h1A5B;
            14'd 9948: out = 14'h1A5A;
            14'd 9949: out = 14'h1A59;
            14'd 9950: out = 14'h1A59;
            14'd 9951: out = 14'h1A58;
            14'd 9952: out = 14'h1A57;
            14'd 9953: out = 14'h1A57;
            14'd 9954: out = 14'h1A56;
            14'd 9955: out = 14'h1A55;
            14'd 9956: out = 14'h1A55;
            14'd 9957: out = 14'h1A54;
            14'd 9958: out = 14'h1A53;
            14'd 9959: out = 14'h1A53;
            14'd 9960: out = 14'h1A52;
            14'd 9961: out = 14'h1A51;
            14'd 9962: out = 14'h1A50;
            14'd 9963: out = 14'h1A50;
            14'd 9964: out = 14'h1A4F;
            14'd 9965: out = 14'h1A4E;
            14'd 9966: out = 14'h1A4E;
            14'd 9967: out = 14'h1A4D;
            14'd 9968: out = 14'h1A4C;
            14'd 9969: out = 14'h1A4C;
            14'd 9970: out = 14'h1A4B;
            14'd 9971: out = 14'h1A4A;
            14'd 9972: out = 14'h1A4A;
            14'd 9973: out = 14'h1A49;
            14'd 9974: out = 14'h1A48;
            14'd 9975: out = 14'h1A48;
            14'd 9976: out = 14'h1A47;
            14'd 9977: out = 14'h1A46;
            14'd 9978: out = 14'h1A46;
            14'd 9979: out = 14'h1A45;
            14'd 9980: out = 14'h1A44;
            14'd 9981: out = 14'h1A44;
            14'd 9982: out = 14'h1A43;
            14'd 9983: out = 14'h1A42;
            14'd 9984: out = 14'h1A42;
            14'd 9985: out = 14'h1A41;
            14'd 9986: out = 14'h1A40;
            14'd 9987: out = 14'h1A40;
            14'd 9988: out = 14'h1A3F;
            14'd 9989: out = 14'h1A3E;
            14'd 9990: out = 14'h1A3E;
            14'd 9991: out = 14'h1A3D;
            14'd 9992: out = 14'h1A3C;
            14'd 9993: out = 14'h1A3C;
            14'd 9994: out = 14'h1A3B;
            14'd 9995: out = 14'h1A3A;
            14'd 9996: out = 14'h1A3A;
            14'd 9997: out = 14'h1A39;
            14'd 9998: out = 14'h1A38;
            14'd 9999: out = 14'h1A38;
            14'd10000: out = 14'h1A37;
            14'd10001: out = 14'h1A36;
            14'd10002: out = 14'h1A36;
            14'd10003: out = 14'h1A35;
            14'd10004: out = 14'h1A34;
            14'd10005: out = 14'h1A34;
            14'd10006: out = 14'h1A33;
            14'd10007: out = 14'h1A32;
            14'd10008: out = 14'h1A32;
            14'd10009: out = 14'h1A31;
            14'd10010: out = 14'h1A30;
            14'd10011: out = 14'h1A30;
            14'd10012: out = 14'h1A2F;
            14'd10013: out = 14'h1A2E;
            14'd10014: out = 14'h1A2E;
            14'd10015: out = 14'h1A2D;
            14'd10016: out = 14'h1A2C;
            14'd10017: out = 14'h1A2B;
            14'd10018: out = 14'h1A2B;
            14'd10019: out = 14'h1A2A;
            14'd10020: out = 14'h1A29;
            14'd10021: out = 14'h1A29;
            14'd10022: out = 14'h1A28;
            14'd10023: out = 14'h1A27;
            14'd10024: out = 14'h1A27;
            14'd10025: out = 14'h1A26;
            14'd10026: out = 14'h1A25;
            14'd10027: out = 14'h1A25;
            14'd10028: out = 14'h1A24;
            14'd10029: out = 14'h1A23;
            14'd10030: out = 14'h1A23;
            14'd10031: out = 14'h1A22;
            14'd10032: out = 14'h1A21;
            14'd10033: out = 14'h1A21;
            14'd10034: out = 14'h1A20;
            14'd10035: out = 14'h1A1F;
            14'd10036: out = 14'h1A1F;
            14'd10037: out = 14'h1A1E;
            14'd10038: out = 14'h1A1D;
            14'd10039: out = 14'h1A1D;
            14'd10040: out = 14'h1A1C;
            14'd10041: out = 14'h1A1B;
            14'd10042: out = 14'h1A1B;
            14'd10043: out = 14'h1A1A;
            14'd10044: out = 14'h1A19;
            14'd10045: out = 14'h1A19;
            14'd10046: out = 14'h1A18;
            14'd10047: out = 14'h1A17;
            14'd10048: out = 14'h1A17;
            14'd10049: out = 14'h1A16;
            14'd10050: out = 14'h1A15;
            14'd10051: out = 14'h1A15;
            14'd10052: out = 14'h1A14;
            14'd10053: out = 14'h1A14;
            14'd10054: out = 14'h1A13;
            14'd10055: out = 14'h1A12;
            14'd10056: out = 14'h1A12;
            14'd10057: out = 14'h1A11;
            14'd10058: out = 14'h1A10;
            14'd10059: out = 14'h1A10;
            14'd10060: out = 14'h1A0F;
            14'd10061: out = 14'h1A0E;
            14'd10062: out = 14'h1A0E;
            14'd10063: out = 14'h1A0D;
            14'd10064: out = 14'h1A0C;
            14'd10065: out = 14'h1A0C;
            14'd10066: out = 14'h1A0B;
            14'd10067: out = 14'h1A0A;
            14'd10068: out = 14'h1A0A;
            14'd10069: out = 14'h1A09;
            14'd10070: out = 14'h1A08;
            14'd10071: out = 14'h1A08;
            14'd10072: out = 14'h1A07;
            14'd10073: out = 14'h1A06;
            14'd10074: out = 14'h1A06;
            14'd10075: out = 14'h1A05;
            14'd10076: out = 14'h1A04;
            14'd10077: out = 14'h1A04;
            14'd10078: out = 14'h1A03;
            14'd10079: out = 14'h1A02;
            14'd10080: out = 14'h1A02;
            14'd10081: out = 14'h1A01;
            14'd10082: out = 14'h1A00;
            14'd10083: out = 14'h1A00;
            14'd10084: out = 14'h19FF;
            14'd10085: out = 14'h19FE;
            14'd10086: out = 14'h19FE;
            14'd10087: out = 14'h19FD;
            14'd10088: out = 14'h19FC;
            14'd10089: out = 14'h19FC;
            14'd10090: out = 14'h19FB;
            14'd10091: out = 14'h19FA;
            14'd10092: out = 14'h19FA;
            14'd10093: out = 14'h19F9;
            14'd10094: out = 14'h19F8;
            14'd10095: out = 14'h19F8;
            14'd10096: out = 14'h19F7;
            14'd10097: out = 14'h19F6;
            14'd10098: out = 14'h19F6;
            14'd10099: out = 14'h19F5;
            14'd10100: out = 14'h19F4;
            14'd10101: out = 14'h19F4;
            14'd10102: out = 14'h19F3;
            14'd10103: out = 14'h19F2;
            14'd10104: out = 14'h19F2;
            14'd10105: out = 14'h19F1;
            14'd10106: out = 14'h19F0;
            14'd10107: out = 14'h19F0;
            14'd10108: out = 14'h19EF;
            14'd10109: out = 14'h19EF;
            14'd10110: out = 14'h19EE;
            14'd10111: out = 14'h19ED;
            14'd10112: out = 14'h19ED;
            14'd10113: out = 14'h19EC;
            14'd10114: out = 14'h19EB;
            14'd10115: out = 14'h19EB;
            14'd10116: out = 14'h19EA;
            14'd10117: out = 14'h19E9;
            14'd10118: out = 14'h19E9;
            14'd10119: out = 14'h19E8;
            14'd10120: out = 14'h19E7;
            14'd10121: out = 14'h19E7;
            14'd10122: out = 14'h19E6;
            14'd10123: out = 14'h19E5;
            14'd10124: out = 14'h19E5;
            14'd10125: out = 14'h19E4;
            14'd10126: out = 14'h19E3;
            14'd10127: out = 14'h19E3;
            14'd10128: out = 14'h19E2;
            14'd10129: out = 14'h19E1;
            14'd10130: out = 14'h19E1;
            14'd10131: out = 14'h19E0;
            14'd10132: out = 14'h19DF;
            14'd10133: out = 14'h19DF;
            14'd10134: out = 14'h19DE;
            14'd10135: out = 14'h19DD;
            14'd10136: out = 14'h19DD;
            14'd10137: out = 14'h19DC;
            14'd10138: out = 14'h19DC;
            14'd10139: out = 14'h19DB;
            14'd10140: out = 14'h19DA;
            14'd10141: out = 14'h19DA;
            14'd10142: out = 14'h19D9;
            14'd10143: out = 14'h19D8;
            14'd10144: out = 14'h19D8;
            14'd10145: out = 14'h19D7;
            14'd10146: out = 14'h19D6;
            14'd10147: out = 14'h19D6;
            14'd10148: out = 14'h19D5;
            14'd10149: out = 14'h19D4;
            14'd10150: out = 14'h19D4;
            14'd10151: out = 14'h19D3;
            14'd10152: out = 14'h19D2;
            14'd10153: out = 14'h19D2;
            14'd10154: out = 14'h19D1;
            14'd10155: out = 14'h19D0;
            14'd10156: out = 14'h19D0;
            14'd10157: out = 14'h19CF;
            14'd10158: out = 14'h19CF;
            14'd10159: out = 14'h19CE;
            14'd10160: out = 14'h19CD;
            14'd10161: out = 14'h19CD;
            14'd10162: out = 14'h19CC;
            14'd10163: out = 14'h19CB;
            14'd10164: out = 14'h19CB;
            14'd10165: out = 14'h19CA;
            14'd10166: out = 14'h19C9;
            14'd10167: out = 14'h19C9;
            14'd10168: out = 14'h19C8;
            14'd10169: out = 14'h19C7;
            14'd10170: out = 14'h19C7;
            14'd10171: out = 14'h19C6;
            14'd10172: out = 14'h19C5;
            14'd10173: out = 14'h19C5;
            14'd10174: out = 14'h19C4;
            14'd10175: out = 14'h19C3;
            14'd10176: out = 14'h19C3;
            14'd10177: out = 14'h19C2;
            14'd10178: out = 14'h19C2;
            14'd10179: out = 14'h19C1;
            14'd10180: out = 14'h19C0;
            14'd10181: out = 14'h19C0;
            14'd10182: out = 14'h19BF;
            14'd10183: out = 14'h19BE;
            14'd10184: out = 14'h19BE;
            14'd10185: out = 14'h19BD;
            14'd10186: out = 14'h19BC;
            14'd10187: out = 14'h19BC;
            14'd10188: out = 14'h19BB;
            14'd10189: out = 14'h19BA;
            14'd10190: out = 14'h19BA;
            14'd10191: out = 14'h19B9;
            14'd10192: out = 14'h19B8;
            14'd10193: out = 14'h19B8;
            14'd10194: out = 14'h19B7;
            14'd10195: out = 14'h19B7;
            14'd10196: out = 14'h19B6;
            14'd10197: out = 14'h19B5;
            14'd10198: out = 14'h19B5;
            14'd10199: out = 14'h19B4;
            14'd10200: out = 14'h19B3;
            14'd10201: out = 14'h19B3;
            14'd10202: out = 14'h19B2;
            14'd10203: out = 14'h19B1;
            14'd10204: out = 14'h19B1;
            14'd10205: out = 14'h19B0;
            14'd10206: out = 14'h19AF;
            14'd10207: out = 14'h19AF;
            14'd10208: out = 14'h19AE;
            14'd10209: out = 14'h19AE;
            14'd10210: out = 14'h19AD;
            14'd10211: out = 14'h19AC;
            14'd10212: out = 14'h19AC;
            14'd10213: out = 14'h19AB;
            14'd10214: out = 14'h19AA;
            14'd10215: out = 14'h19AA;
            14'd10216: out = 14'h19A9;
            14'd10217: out = 14'h19A8;
            14'd10218: out = 14'h19A8;
            14'd10219: out = 14'h19A7;
            14'd10220: out = 14'h19A6;
            14'd10221: out = 14'h19A6;
            14'd10222: out = 14'h19A5;
            14'd10223: out = 14'h19A4;
            14'd10224: out = 14'h19A4;
            14'd10225: out = 14'h19A3;
            14'd10226: out = 14'h19A3;
            14'd10227: out = 14'h19A2;
            14'd10228: out = 14'h19A1;
            14'd10229: out = 14'h19A1;
            14'd10230: out = 14'h19A0;
            14'd10231: out = 14'h199F;
            14'd10232: out = 14'h199F;
            14'd10233: out = 14'h199E;
            14'd10234: out = 14'h199D;
            14'd10235: out = 14'h199D;
            14'd10236: out = 14'h199C;
            14'd10237: out = 14'h199C;
            14'd10238: out = 14'h199B;
            14'd10239: out = 14'h199A;
            14'd10240: out = 14'h199A;
            14'd10241: out = 14'h1999;
            14'd10242: out = 14'h1998;
            14'd10243: out = 14'h1998;
            14'd10244: out = 14'h1997;
            14'd10245: out = 14'h1996;
            14'd10246: out = 14'h1996;
            14'd10247: out = 14'h1995;
            14'd10248: out = 14'h1994;
            14'd10249: out = 14'h1994;
            14'd10250: out = 14'h1993;
            14'd10251: out = 14'h1993;
            14'd10252: out = 14'h1992;
            14'd10253: out = 14'h1991;
            14'd10254: out = 14'h1991;
            14'd10255: out = 14'h1990;
            14'd10256: out = 14'h198F;
            14'd10257: out = 14'h198F;
            14'd10258: out = 14'h198E;
            14'd10259: out = 14'h198D;
            14'd10260: out = 14'h198D;
            14'd10261: out = 14'h198C;
            14'd10262: out = 14'h198C;
            14'd10263: out = 14'h198B;
            14'd10264: out = 14'h198A;
            14'd10265: out = 14'h198A;
            14'd10266: out = 14'h1989;
            14'd10267: out = 14'h1988;
            14'd10268: out = 14'h1988;
            14'd10269: out = 14'h1987;
            14'd10270: out = 14'h1986;
            14'd10271: out = 14'h1986;
            14'd10272: out = 14'h1985;
            14'd10273: out = 14'h1985;
            14'd10274: out = 14'h1984;
            14'd10275: out = 14'h1983;
            14'd10276: out = 14'h1983;
            14'd10277: out = 14'h1982;
            14'd10278: out = 14'h1981;
            14'd10279: out = 14'h1981;
            14'd10280: out = 14'h1980;
            14'd10281: out = 14'h197F;
            14'd10282: out = 14'h197F;
            14'd10283: out = 14'h197E;
            14'd10284: out = 14'h197E;
            14'd10285: out = 14'h197D;
            14'd10286: out = 14'h197C;
            14'd10287: out = 14'h197C;
            14'd10288: out = 14'h197B;
            14'd10289: out = 14'h197A;
            14'd10290: out = 14'h197A;
            14'd10291: out = 14'h1979;
            14'd10292: out = 14'h1978;
            14'd10293: out = 14'h1978;
            14'd10294: out = 14'h1977;
            14'd10295: out = 14'h1977;
            14'd10296: out = 14'h1976;
            14'd10297: out = 14'h1975;
            14'd10298: out = 14'h1975;
            14'd10299: out = 14'h1974;
            14'd10300: out = 14'h1973;
            14'd10301: out = 14'h1973;
            14'd10302: out = 14'h1972;
            14'd10303: out = 14'h1972;
            14'd10304: out = 14'h1971;
            14'd10305: out = 14'h1970;
            14'd10306: out = 14'h1970;
            14'd10307: out = 14'h196F;
            14'd10308: out = 14'h196E;
            14'd10309: out = 14'h196E;
            14'd10310: out = 14'h196D;
            14'd10311: out = 14'h196C;
            14'd10312: out = 14'h196C;
            14'd10313: out = 14'h196B;
            14'd10314: out = 14'h196B;
            14'd10315: out = 14'h196A;
            14'd10316: out = 14'h1969;
            14'd10317: out = 14'h1969;
            14'd10318: out = 14'h1968;
            14'd10319: out = 14'h1967;
            14'd10320: out = 14'h1967;
            14'd10321: out = 14'h1966;
            14'd10322: out = 14'h1966;
            14'd10323: out = 14'h1965;
            14'd10324: out = 14'h1964;
            14'd10325: out = 14'h1964;
            14'd10326: out = 14'h1963;
            14'd10327: out = 14'h1962;
            14'd10328: out = 14'h1962;
            14'd10329: out = 14'h1961;
            14'd10330: out = 14'h1961;
            14'd10331: out = 14'h1960;
            14'd10332: out = 14'h195F;
            14'd10333: out = 14'h195F;
            14'd10334: out = 14'h195E;
            14'd10335: out = 14'h195D;
            14'd10336: out = 14'h195D;
            14'd10337: out = 14'h195C;
            14'd10338: out = 14'h195B;
            14'd10339: out = 14'h195B;
            14'd10340: out = 14'h195A;
            14'd10341: out = 14'h195A;
            14'd10342: out = 14'h1959;
            14'd10343: out = 14'h1958;
            14'd10344: out = 14'h1958;
            14'd10345: out = 14'h1957;
            14'd10346: out = 14'h1956;
            14'd10347: out = 14'h1956;
            14'd10348: out = 14'h1955;
            14'd10349: out = 14'h1955;
            14'd10350: out = 14'h1954;
            14'd10351: out = 14'h1953;
            14'd10352: out = 14'h1953;
            14'd10353: out = 14'h1952;
            14'd10354: out = 14'h1951;
            14'd10355: out = 14'h1951;
            14'd10356: out = 14'h1950;
            14'd10357: out = 14'h1950;
            14'd10358: out = 14'h194F;
            14'd10359: out = 14'h194E;
            14'd10360: out = 14'h194E;
            14'd10361: out = 14'h194D;
            14'd10362: out = 14'h194C;
            14'd10363: out = 14'h194C;
            14'd10364: out = 14'h194B;
            14'd10365: out = 14'h194B;
            14'd10366: out = 14'h194A;
            14'd10367: out = 14'h1949;
            14'd10368: out = 14'h1949;
            14'd10369: out = 14'h1948;
            14'd10370: out = 14'h1947;
            14'd10371: out = 14'h1947;
            14'd10372: out = 14'h1946;
            14'd10373: out = 14'h1946;
            14'd10374: out = 14'h1945;
            14'd10375: out = 14'h1944;
            14'd10376: out = 14'h1944;
            14'd10377: out = 14'h1943;
            14'd10378: out = 14'h1942;
            14'd10379: out = 14'h1942;
            14'd10380: out = 14'h1941;
            14'd10381: out = 14'h1941;
            14'd10382: out = 14'h1940;
            14'd10383: out = 14'h193F;
            14'd10384: out = 14'h193F;
            14'd10385: out = 14'h193E;
            14'd10386: out = 14'h193D;
            14'd10387: out = 14'h193D;
            14'd10388: out = 14'h193C;
            14'd10389: out = 14'h193C;
            14'd10390: out = 14'h193B;
            14'd10391: out = 14'h193A;
            14'd10392: out = 14'h193A;
            14'd10393: out = 14'h1939;
            14'd10394: out = 14'h1939;
            14'd10395: out = 14'h1938;
            14'd10396: out = 14'h1937;
            14'd10397: out = 14'h1937;
            14'd10398: out = 14'h1936;
            14'd10399: out = 14'h1935;
            14'd10400: out = 14'h1935;
            14'd10401: out = 14'h1934;
            14'd10402: out = 14'h1934;
            14'd10403: out = 14'h1933;
            14'd10404: out = 14'h1932;
            14'd10405: out = 14'h1932;
            14'd10406: out = 14'h1931;
            14'd10407: out = 14'h1930;
            14'd10408: out = 14'h1930;
            14'd10409: out = 14'h192F;
            14'd10410: out = 14'h192F;
            14'd10411: out = 14'h192E;
            14'd10412: out = 14'h192D;
            14'd10413: out = 14'h192D;
            14'd10414: out = 14'h192C;
            14'd10415: out = 14'h192B;
            14'd10416: out = 14'h192B;
            14'd10417: out = 14'h192A;
            14'd10418: out = 14'h192A;
            14'd10419: out = 14'h1929;
            14'd10420: out = 14'h1928;
            14'd10421: out = 14'h1928;
            14'd10422: out = 14'h1927;
            14'd10423: out = 14'h1927;
            14'd10424: out = 14'h1926;
            14'd10425: out = 14'h1925;
            14'd10426: out = 14'h1925;
            14'd10427: out = 14'h1924;
            14'd10428: out = 14'h1923;
            14'd10429: out = 14'h1923;
            14'd10430: out = 14'h1922;
            14'd10431: out = 14'h1922;
            14'd10432: out = 14'h1921;
            14'd10433: out = 14'h1920;
            14'd10434: out = 14'h1920;
            14'd10435: out = 14'h191F;
            14'd10436: out = 14'h191F;
            14'd10437: out = 14'h191E;
            14'd10438: out = 14'h191D;
            14'd10439: out = 14'h191D;
            14'd10440: out = 14'h191C;
            14'd10441: out = 14'h191B;
            14'd10442: out = 14'h191B;
            14'd10443: out = 14'h191A;
            14'd10444: out = 14'h191A;
            14'd10445: out = 14'h1919;
            14'd10446: out = 14'h1918;
            14'd10447: out = 14'h1918;
            14'd10448: out = 14'h1917;
            14'd10449: out = 14'h1917;
            14'd10450: out = 14'h1916;
            14'd10451: out = 14'h1915;
            14'd10452: out = 14'h1915;
            14'd10453: out = 14'h1914;
            14'd10454: out = 14'h1913;
            14'd10455: out = 14'h1913;
            14'd10456: out = 14'h1912;
            14'd10457: out = 14'h1912;
            14'd10458: out = 14'h1911;
            14'd10459: out = 14'h1910;
            14'd10460: out = 14'h1910;
            14'd10461: out = 14'h190F;
            14'd10462: out = 14'h190F;
            14'd10463: out = 14'h190E;
            14'd10464: out = 14'h190D;
            14'd10465: out = 14'h190D;
            14'd10466: out = 14'h190C;
            14'd10467: out = 14'h190B;
            14'd10468: out = 14'h190B;
            14'd10469: out = 14'h190A;
            14'd10470: out = 14'h190A;
            14'd10471: out = 14'h1909;
            14'd10472: out = 14'h1908;
            14'd10473: out = 14'h1908;
            14'd10474: out = 14'h1907;
            14'd10475: out = 14'h1907;
            14'd10476: out = 14'h1906;
            14'd10477: out = 14'h1905;
            14'd10478: out = 14'h1905;
            14'd10479: out = 14'h1904;
            14'd10480: out = 14'h1904;
            14'd10481: out = 14'h1903;
            14'd10482: out = 14'h1902;
            14'd10483: out = 14'h1902;
            14'd10484: out = 14'h1901;
            14'd10485: out = 14'h1900;
            14'd10486: out = 14'h1900;
            14'd10487: out = 14'h18FF;
            14'd10488: out = 14'h18FF;
            14'd10489: out = 14'h18FE;
            14'd10490: out = 14'h18FD;
            14'd10491: out = 14'h18FD;
            14'd10492: out = 14'h18FC;
            14'd10493: out = 14'h18FC;
            14'd10494: out = 14'h18FB;
            14'd10495: out = 14'h18FA;
            14'd10496: out = 14'h18FA;
            14'd10497: out = 14'h18F9;
            14'd10498: out = 14'h18F9;
            14'd10499: out = 14'h18F8;
            14'd10500: out = 14'h18F7;
            14'd10501: out = 14'h18F7;
            14'd10502: out = 14'h18F6;
            14'd10503: out = 14'h18F5;
            14'd10504: out = 14'h18F5;
            14'd10505: out = 14'h18F4;
            14'd10506: out = 14'h18F4;
            14'd10507: out = 14'h18F3;
            14'd10508: out = 14'h18F2;
            14'd10509: out = 14'h18F2;
            14'd10510: out = 14'h18F1;
            14'd10511: out = 14'h18F1;
            14'd10512: out = 14'h18F0;
            14'd10513: out = 14'h18EF;
            14'd10514: out = 14'h18EF;
            14'd10515: out = 14'h18EE;
            14'd10516: out = 14'h18EE;
            14'd10517: out = 14'h18ED;
            14'd10518: out = 14'h18EC;
            14'd10519: out = 14'h18EC;
            14'd10520: out = 14'h18EB;
            14'd10521: out = 14'h18EB;
            14'd10522: out = 14'h18EA;
            14'd10523: out = 14'h18E9;
            14'd10524: out = 14'h18E9;
            14'd10525: out = 14'h18E8;
            14'd10526: out = 14'h18E8;
            14'd10527: out = 14'h18E7;
            14'd10528: out = 14'h18E6;
            14'd10529: out = 14'h18E6;
            14'd10530: out = 14'h18E5;
            14'd10531: out = 14'h18E5;
            14'd10532: out = 14'h18E4;
            14'd10533: out = 14'h18E3;
            14'd10534: out = 14'h18E3;
            14'd10535: out = 14'h18E2;
            14'd10536: out = 14'h18E1;
            14'd10537: out = 14'h18E1;
            14'd10538: out = 14'h18E0;
            14'd10539: out = 14'h18E0;
            14'd10540: out = 14'h18DF;
            14'd10541: out = 14'h18DE;
            14'd10542: out = 14'h18DE;
            14'd10543: out = 14'h18DD;
            14'd10544: out = 14'h18DD;
            14'd10545: out = 14'h18DC;
            14'd10546: out = 14'h18DB;
            14'd10547: out = 14'h18DB;
            14'd10548: out = 14'h18DA;
            14'd10549: out = 14'h18DA;
            14'd10550: out = 14'h18D9;
            14'd10551: out = 14'h18D8;
            14'd10552: out = 14'h18D8;
            14'd10553: out = 14'h18D7;
            14'd10554: out = 14'h18D7;
            14'd10555: out = 14'h18D6;
            14'd10556: out = 14'h18D5;
            14'd10557: out = 14'h18D5;
            14'd10558: out = 14'h18D4;
            14'd10559: out = 14'h18D4;
            14'd10560: out = 14'h18D3;
            14'd10561: out = 14'h18D2;
            14'd10562: out = 14'h18D2;
            14'd10563: out = 14'h18D1;
            14'd10564: out = 14'h18D1;
            14'd10565: out = 14'h18D0;
            14'd10566: out = 14'h18CF;
            14'd10567: out = 14'h18CF;
            14'd10568: out = 14'h18CE;
            14'd10569: out = 14'h18CE;
            14'd10570: out = 14'h18CD;
            14'd10571: out = 14'h18CC;
            14'd10572: out = 14'h18CC;
            14'd10573: out = 14'h18CB;
            14'd10574: out = 14'h18CB;
            14'd10575: out = 14'h18CA;
            14'd10576: out = 14'h18C9;
            14'd10577: out = 14'h18C9;
            14'd10578: out = 14'h18C8;
            14'd10579: out = 14'h18C8;
            14'd10580: out = 14'h18C7;
            14'd10581: out = 14'h18C6;
            14'd10582: out = 14'h18C6;
            14'd10583: out = 14'h18C5;
            14'd10584: out = 14'h18C5;
            14'd10585: out = 14'h18C4;
            14'd10586: out = 14'h18C3;
            14'd10587: out = 14'h18C3;
            14'd10588: out = 14'h18C2;
            14'd10589: out = 14'h18C2;
            14'd10590: out = 14'h18C1;
            14'd10591: out = 14'h18C0;
            14'd10592: out = 14'h18C0;
            14'd10593: out = 14'h18BF;
            14'd10594: out = 14'h18BF;
            14'd10595: out = 14'h18BE;
            14'd10596: out = 14'h18BD;
            14'd10597: out = 14'h18BD;
            14'd10598: out = 14'h18BC;
            14'd10599: out = 14'h18BC;
            14'd10600: out = 14'h18BB;
            14'd10601: out = 14'h18BA;
            14'd10602: out = 14'h18BA;
            14'd10603: out = 14'h18B9;
            14'd10604: out = 14'h18B9;
            14'd10605: out = 14'h18B8;
            14'd10606: out = 14'h18B7;
            14'd10607: out = 14'h18B7;
            14'd10608: out = 14'h18B6;
            14'd10609: out = 14'h18B6;
            14'd10610: out = 14'h18B5;
            14'd10611: out = 14'h18B4;
            14'd10612: out = 14'h18B4;
            14'd10613: out = 14'h18B3;
            14'd10614: out = 14'h18B3;
            14'd10615: out = 14'h18B2;
            14'd10616: out = 14'h18B1;
            14'd10617: out = 14'h18B1;
            14'd10618: out = 14'h18B0;
            14'd10619: out = 14'h18B0;
            14'd10620: out = 14'h18AF;
            14'd10621: out = 14'h18AF;
            14'd10622: out = 14'h18AE;
            14'd10623: out = 14'h18AD;
            14'd10624: out = 14'h18AD;
            14'd10625: out = 14'h18AC;
            14'd10626: out = 14'h18AC;
            14'd10627: out = 14'h18AB;
            14'd10628: out = 14'h18AA;
            14'd10629: out = 14'h18AA;
            14'd10630: out = 14'h18A9;
            14'd10631: out = 14'h18A9;
            14'd10632: out = 14'h18A8;
            14'd10633: out = 14'h18A7;
            14'd10634: out = 14'h18A7;
            14'd10635: out = 14'h18A6;
            14'd10636: out = 14'h18A6;
            14'd10637: out = 14'h18A5;
            14'd10638: out = 14'h18A4;
            14'd10639: out = 14'h18A4;
            14'd10640: out = 14'h18A3;
            14'd10641: out = 14'h18A3;
            14'd10642: out = 14'h18A2;
            14'd10643: out = 14'h18A1;
            14'd10644: out = 14'h18A1;
            14'd10645: out = 14'h18A0;
            14'd10646: out = 14'h18A0;
            14'd10647: out = 14'h189F;
            14'd10648: out = 14'h189E;
            14'd10649: out = 14'h189E;
            14'd10650: out = 14'h189D;
            14'd10651: out = 14'h189D;
            14'd10652: out = 14'h189C;
            14'd10653: out = 14'h189C;
            14'd10654: out = 14'h189B;
            14'd10655: out = 14'h189A;
            14'd10656: out = 14'h189A;
            14'd10657: out = 14'h1899;
            14'd10658: out = 14'h1899;
            14'd10659: out = 14'h1898;
            14'd10660: out = 14'h1897;
            14'd10661: out = 14'h1897;
            14'd10662: out = 14'h1896;
            14'd10663: out = 14'h1896;
            14'd10664: out = 14'h1895;
            14'd10665: out = 14'h1894;
            14'd10666: out = 14'h1894;
            14'd10667: out = 14'h1893;
            14'd10668: out = 14'h1893;
            14'd10669: out = 14'h1892;
            14'd10670: out = 14'h1891;
            14'd10671: out = 14'h1891;
            14'd10672: out = 14'h1890;
            14'd10673: out = 14'h1890;
            14'd10674: out = 14'h188F;
            14'd10675: out = 14'h188F;
            14'd10676: out = 14'h188E;
            14'd10677: out = 14'h188D;
            14'd10678: out = 14'h188D;
            14'd10679: out = 14'h188C;
            14'd10680: out = 14'h188C;
            14'd10681: out = 14'h188B;
            14'd10682: out = 14'h188A;
            14'd10683: out = 14'h188A;
            14'd10684: out = 14'h1889;
            14'd10685: out = 14'h1889;
            14'd10686: out = 14'h1888;
            14'd10687: out = 14'h1887;
            14'd10688: out = 14'h1887;
            14'd10689: out = 14'h1886;
            14'd10690: out = 14'h1886;
            14'd10691: out = 14'h1885;
            14'd10692: out = 14'h1885;
            14'd10693: out = 14'h1884;
            14'd10694: out = 14'h1883;
            14'd10695: out = 14'h1883;
            14'd10696: out = 14'h1882;
            14'd10697: out = 14'h1882;
            14'd10698: out = 14'h1881;
            14'd10699: out = 14'h1880;
            14'd10700: out = 14'h1880;
            14'd10701: out = 14'h187F;
            14'd10702: out = 14'h187F;
            14'd10703: out = 14'h187E;
            14'd10704: out = 14'h187E;
            14'd10705: out = 14'h187D;
            14'd10706: out = 14'h187C;
            14'd10707: out = 14'h187C;
            14'd10708: out = 14'h187B;
            14'd10709: out = 14'h187B;
            14'd10710: out = 14'h187A;
            14'd10711: out = 14'h1879;
            14'd10712: out = 14'h1879;
            14'd10713: out = 14'h1878;
            14'd10714: out = 14'h1878;
            14'd10715: out = 14'h1877;
            14'd10716: out = 14'h1876;
            14'd10717: out = 14'h1876;
            14'd10718: out = 14'h1875;
            14'd10719: out = 14'h1875;
            14'd10720: out = 14'h1874;
            14'd10721: out = 14'h1874;
            14'd10722: out = 14'h1873;
            14'd10723: out = 14'h1872;
            14'd10724: out = 14'h1872;
            14'd10725: out = 14'h1871;
            14'd10726: out = 14'h1871;
            14'd10727: out = 14'h1870;
            14'd10728: out = 14'h186F;
            14'd10729: out = 14'h186F;
            14'd10730: out = 14'h186E;
            14'd10731: out = 14'h186E;
            14'd10732: out = 14'h186D;
            14'd10733: out = 14'h186D;
            14'd10734: out = 14'h186C;
            14'd10735: out = 14'h186B;
            14'd10736: out = 14'h186B;
            14'd10737: out = 14'h186A;
            14'd10738: out = 14'h186A;
            14'd10739: out = 14'h1869;
            14'd10740: out = 14'h1868;
            14'd10741: out = 14'h1868;
            14'd10742: out = 14'h1867;
            14'd10743: out = 14'h1867;
            14'd10744: out = 14'h1866;
            14'd10745: out = 14'h1866;
            14'd10746: out = 14'h1865;
            14'd10747: out = 14'h1864;
            14'd10748: out = 14'h1864;
            14'd10749: out = 14'h1863;
            14'd10750: out = 14'h1863;
            14'd10751: out = 14'h1862;
            14'd10752: out = 14'h1862;
            14'd10753: out = 14'h1861;
            14'd10754: out = 14'h1860;
            14'd10755: out = 14'h1860;
            14'd10756: out = 14'h185F;
            14'd10757: out = 14'h185F;
            14'd10758: out = 14'h185E;
            14'd10759: out = 14'h185D;
            14'd10760: out = 14'h185D;
            14'd10761: out = 14'h185C;
            14'd10762: out = 14'h185C;
            14'd10763: out = 14'h185B;
            14'd10764: out = 14'h185B;
            14'd10765: out = 14'h185A;
            14'd10766: out = 14'h1859;
            14'd10767: out = 14'h1859;
            14'd10768: out = 14'h1858;
            14'd10769: out = 14'h1858;
            14'd10770: out = 14'h1857;
            14'd10771: out = 14'h1857;
            14'd10772: out = 14'h1856;
            14'd10773: out = 14'h1855;
            14'd10774: out = 14'h1855;
            14'd10775: out = 14'h1854;
            14'd10776: out = 14'h1854;
            14'd10777: out = 14'h1853;
            14'd10778: out = 14'h1852;
            14'd10779: out = 14'h1852;
            14'd10780: out = 14'h1851;
            14'd10781: out = 14'h1851;
            14'd10782: out = 14'h1850;
            14'd10783: out = 14'h1850;
            14'd10784: out = 14'h184F;
            14'd10785: out = 14'h184E;
            14'd10786: out = 14'h184E;
            14'd10787: out = 14'h184D;
            14'd10788: out = 14'h184D;
            14'd10789: out = 14'h184C;
            14'd10790: out = 14'h184C;
            14'd10791: out = 14'h184B;
            14'd10792: out = 14'h184A;
            14'd10793: out = 14'h184A;
            14'd10794: out = 14'h1849;
            14'd10795: out = 14'h1849;
            14'd10796: out = 14'h1848;
            14'd10797: out = 14'h1848;
            14'd10798: out = 14'h1847;
            14'd10799: out = 14'h1846;
            14'd10800: out = 14'h1846;
            14'd10801: out = 14'h1845;
            14'd10802: out = 14'h1845;
            14'd10803: out = 14'h1844;
            14'd10804: out = 14'h1843;
            14'd10805: out = 14'h1843;
            14'd10806: out = 14'h1842;
            14'd10807: out = 14'h1842;
            14'd10808: out = 14'h1841;
            14'd10809: out = 14'h1841;
            14'd10810: out = 14'h1840;
            14'd10811: out = 14'h183F;
            14'd10812: out = 14'h183F;
            14'd10813: out = 14'h183E;
            14'd10814: out = 14'h183E;
            14'd10815: out = 14'h183D;
            14'd10816: out = 14'h183D;
            14'd10817: out = 14'h183C;
            14'd10818: out = 14'h183B;
            14'd10819: out = 14'h183B;
            14'd10820: out = 14'h183A;
            14'd10821: out = 14'h183A;
            14'd10822: out = 14'h1839;
            14'd10823: out = 14'h1839;
            14'd10824: out = 14'h1838;
            14'd10825: out = 14'h1837;
            14'd10826: out = 14'h1837;
            14'd10827: out = 14'h1836;
            14'd10828: out = 14'h1836;
            14'd10829: out = 14'h1835;
            14'd10830: out = 14'h1835;
            14'd10831: out = 14'h1834;
            14'd10832: out = 14'h1833;
            14'd10833: out = 14'h1833;
            14'd10834: out = 14'h1832;
            14'd10835: out = 14'h1832;
            14'd10836: out = 14'h1831;
            14'd10837: out = 14'h1831;
            14'd10838: out = 14'h1830;
            14'd10839: out = 14'h182F;
            14'd10840: out = 14'h182F;
            14'd10841: out = 14'h182E;
            14'd10842: out = 14'h182E;
            14'd10843: out = 14'h182D;
            14'd10844: out = 14'h182D;
            14'd10845: out = 14'h182C;
            14'd10846: out = 14'h182B;
            14'd10847: out = 14'h182B;
            14'd10848: out = 14'h182A;
            14'd10849: out = 14'h182A;
            14'd10850: out = 14'h1829;
            14'd10851: out = 14'h1829;
            14'd10852: out = 14'h1828;
            14'd10853: out = 14'h1827;
            14'd10854: out = 14'h1827;
            14'd10855: out = 14'h1826;
            14'd10856: out = 14'h1826;
            14'd10857: out = 14'h1825;
            14'd10858: out = 14'h1825;
            14'd10859: out = 14'h1824;
            14'd10860: out = 14'h1823;
            14'd10861: out = 14'h1823;
            14'd10862: out = 14'h1822;
            14'd10863: out = 14'h1822;
            14'd10864: out = 14'h1821;
            14'd10865: out = 14'h1821;
            14'd10866: out = 14'h1820;
            14'd10867: out = 14'h181F;
            14'd10868: out = 14'h181F;
            14'd10869: out = 14'h181E;
            14'd10870: out = 14'h181E;
            14'd10871: out = 14'h181D;
            14'd10872: out = 14'h181D;
            14'd10873: out = 14'h181C;
            14'd10874: out = 14'h181B;
            14'd10875: out = 14'h181B;
            14'd10876: out = 14'h181A;
            14'd10877: out = 14'h181A;
            14'd10878: out = 14'h1819;
            14'd10879: out = 14'h1819;
            14'd10880: out = 14'h1818;
            14'd10881: out = 14'h1818;
            14'd10882: out = 14'h1817;
            14'd10883: out = 14'h1816;
            14'd10884: out = 14'h1816;
            14'd10885: out = 14'h1815;
            14'd10886: out = 14'h1815;
            14'd10887: out = 14'h1814;
            14'd10888: out = 14'h1814;
            14'd10889: out = 14'h1813;
            14'd10890: out = 14'h1812;
            14'd10891: out = 14'h1812;
            14'd10892: out = 14'h1811;
            14'd10893: out = 14'h1811;
            14'd10894: out = 14'h1810;
            14'd10895: out = 14'h1810;
            14'd10896: out = 14'h180F;
            14'd10897: out = 14'h180E;
            14'd10898: out = 14'h180E;
            14'd10899: out = 14'h180D;
            14'd10900: out = 14'h180D;
            14'd10901: out = 14'h180C;
            14'd10902: out = 14'h180C;
            14'd10903: out = 14'h180B;
            14'd10904: out = 14'h180B;
            14'd10905: out = 14'h180A;
            14'd10906: out = 14'h1809;
            14'd10907: out = 14'h1809;
            14'd10908: out = 14'h1808;
            14'd10909: out = 14'h1808;
            14'd10910: out = 14'h1807;
            14'd10911: out = 14'h1807;
            14'd10912: out = 14'h1806;
            14'd10913: out = 14'h1805;
            14'd10914: out = 14'h1805;
            14'd10915: out = 14'h1804;
            14'd10916: out = 14'h1804;
            14'd10917: out = 14'h1803;
            14'd10918: out = 14'h1803;
            14'd10919: out = 14'h1802;
            14'd10920: out = 14'h1802;
            14'd10921: out = 14'h1801;
            14'd10922: out = 14'h1800;
            14'd10923: out = 14'h1800;
            14'd10924: out = 14'h17FF;
            14'd10925: out = 14'h17FF;
            14'd10926: out = 14'h17FE;
            14'd10927: out = 14'h17FE;
            14'd10928: out = 14'h17FD;
            14'd10929: out = 14'h17FC;
            14'd10930: out = 14'h17FC;
            14'd10931: out = 14'h17FB;
            14'd10932: out = 14'h17FB;
            14'd10933: out = 14'h17FA;
            14'd10934: out = 14'h17FA;
            14'd10935: out = 14'h17F9;
            14'd10936: out = 14'h17F9;
            14'd10937: out = 14'h17F8;
            14'd10938: out = 14'h17F7;
            14'd10939: out = 14'h17F7;
            14'd10940: out = 14'h17F6;
            14'd10941: out = 14'h17F6;
            14'd10942: out = 14'h17F5;
            14'd10943: out = 14'h17F5;
            14'd10944: out = 14'h17F4;
            14'd10945: out = 14'h17F3;
            14'd10946: out = 14'h17F3;
            14'd10947: out = 14'h17F2;
            14'd10948: out = 14'h17F2;
            14'd10949: out = 14'h17F1;
            14'd10950: out = 14'h17F1;
            14'd10951: out = 14'h17F0;
            14'd10952: out = 14'h17F0;
            14'd10953: out = 14'h17EF;
            14'd10954: out = 14'h17EE;
            14'd10955: out = 14'h17EE;
            14'd10956: out = 14'h17ED;
            14'd10957: out = 14'h17ED;
            14'd10958: out = 14'h17EC;
            14'd10959: out = 14'h17EC;
            14'd10960: out = 14'h17EB;
            14'd10961: out = 14'h17EB;
            14'd10962: out = 14'h17EA;
            14'd10963: out = 14'h17E9;
            14'd10964: out = 14'h17E9;
            14'd10965: out = 14'h17E8;
            14'd10966: out = 14'h17E8;
            14'd10967: out = 14'h17E7;
            14'd10968: out = 14'h17E7;
            14'd10969: out = 14'h17E6;
            14'd10970: out = 14'h17E5;
            14'd10971: out = 14'h17E5;
            14'd10972: out = 14'h17E4;
            14'd10973: out = 14'h17E4;
            14'd10974: out = 14'h17E3;
            14'd10975: out = 14'h17E3;
            14'd10976: out = 14'h17E2;
            14'd10977: out = 14'h17E2;
            14'd10978: out = 14'h17E1;
            14'd10979: out = 14'h17E0;
            14'd10980: out = 14'h17E0;
            14'd10981: out = 14'h17DF;
            14'd10982: out = 14'h17DF;
            14'd10983: out = 14'h17DE;
            14'd10984: out = 14'h17DE;
            14'd10985: out = 14'h17DD;
            14'd10986: out = 14'h17DD;
            14'd10987: out = 14'h17DC;
            14'd10988: out = 14'h17DB;
            14'd10989: out = 14'h17DB;
            14'd10990: out = 14'h17DA;
            14'd10991: out = 14'h17DA;
            14'd10992: out = 14'h17D9;
            14'd10993: out = 14'h17D9;
            14'd10994: out = 14'h17D8;
            14'd10995: out = 14'h17D8;
            14'd10996: out = 14'h17D7;
            14'd10997: out = 14'h17D6;
            14'd10998: out = 14'h17D6;
            14'd10999: out = 14'h17D5;
            14'd11000: out = 14'h17D5;
            14'd11001: out = 14'h17D4;
            14'd11002: out = 14'h17D4;
            14'd11003: out = 14'h17D3;
            14'd11004: out = 14'h17D3;
            14'd11005: out = 14'h17D2;
            14'd11006: out = 14'h17D1;
            14'd11007: out = 14'h17D1;
            14'd11008: out = 14'h17D0;
            14'd11009: out = 14'h17D0;
            14'd11010: out = 14'h17CF;
            14'd11011: out = 14'h17CF;
            14'd11012: out = 14'h17CE;
            14'd11013: out = 14'h17CE;
            14'd11014: out = 14'h17CD;
            14'd11015: out = 14'h17CC;
            14'd11016: out = 14'h17CC;
            14'd11017: out = 14'h17CB;
            14'd11018: out = 14'h17CB;
            14'd11019: out = 14'h17CA;
            14'd11020: out = 14'h17CA;
            14'd11021: out = 14'h17C9;
            14'd11022: out = 14'h17C9;
            14'd11023: out = 14'h17C8;
            14'd11024: out = 14'h17C8;
            14'd11025: out = 14'h17C7;
            14'd11026: out = 14'h17C6;
            14'd11027: out = 14'h17C6;
            14'd11028: out = 14'h17C5;
            14'd11029: out = 14'h17C5;
            14'd11030: out = 14'h17C4;
            14'd11031: out = 14'h17C4;
            14'd11032: out = 14'h17C3;
            14'd11033: out = 14'h17C3;
            14'd11034: out = 14'h17C2;
            14'd11035: out = 14'h17C1;
            14'd11036: out = 14'h17C1;
            14'd11037: out = 14'h17C0;
            14'd11038: out = 14'h17C0;
            14'd11039: out = 14'h17BF;
            14'd11040: out = 14'h17BF;
            14'd11041: out = 14'h17BE;
            14'd11042: out = 14'h17BE;
            14'd11043: out = 14'h17BD;
            14'd11044: out = 14'h17BC;
            14'd11045: out = 14'h17BC;
            14'd11046: out = 14'h17BB;
            14'd11047: out = 14'h17BB;
            14'd11048: out = 14'h17BA;
            14'd11049: out = 14'h17BA;
            14'd11050: out = 14'h17B9;
            14'd11051: out = 14'h17B9;
            14'd11052: out = 14'h17B8;
            14'd11053: out = 14'h17B8;
            14'd11054: out = 14'h17B7;
            14'd11055: out = 14'h17B6;
            14'd11056: out = 14'h17B6;
            14'd11057: out = 14'h17B5;
            14'd11058: out = 14'h17B5;
            14'd11059: out = 14'h17B4;
            14'd11060: out = 14'h17B4;
            14'd11061: out = 14'h17B3;
            14'd11062: out = 14'h17B3;
            14'd11063: out = 14'h17B2;
            14'd11064: out = 14'h17B2;
            14'd11065: out = 14'h17B1;
            14'd11066: out = 14'h17B0;
            14'd11067: out = 14'h17B0;
            14'd11068: out = 14'h17AF;
            14'd11069: out = 14'h17AF;
            14'd11070: out = 14'h17AE;
            14'd11071: out = 14'h17AE;
            14'd11072: out = 14'h17AD;
            14'd11073: out = 14'h17AD;
            14'd11074: out = 14'h17AC;
            14'd11075: out = 14'h17AB;
            14'd11076: out = 14'h17AB;
            14'd11077: out = 14'h17AA;
            14'd11078: out = 14'h17AA;
            14'd11079: out = 14'h17A9;
            14'd11080: out = 14'h17A9;
            14'd11081: out = 14'h17A8;
            14'd11082: out = 14'h17A8;
            14'd11083: out = 14'h17A7;
            14'd11084: out = 14'h17A7;
            14'd11085: out = 14'h17A6;
            14'd11086: out = 14'h17A5;
            14'd11087: out = 14'h17A5;
            14'd11088: out = 14'h17A4;
            14'd11089: out = 14'h17A4;
            14'd11090: out = 14'h17A3;
            14'd11091: out = 14'h17A3;
            14'd11092: out = 14'h17A2;
            14'd11093: out = 14'h17A2;
            14'd11094: out = 14'h17A1;
            14'd11095: out = 14'h17A1;
            14'd11096: out = 14'h17A0;
            14'd11097: out = 14'h179F;
            14'd11098: out = 14'h179F;
            14'd11099: out = 14'h179E;
            14'd11100: out = 14'h179E;
            14'd11101: out = 14'h179D;
            14'd11102: out = 14'h179D;
            14'd11103: out = 14'h179C;
            14'd11104: out = 14'h179C;
            14'd11105: out = 14'h179B;
            14'd11106: out = 14'h179B;
            14'd11107: out = 14'h179A;
            14'd11108: out = 14'h1799;
            14'd11109: out = 14'h1799;
            14'd11110: out = 14'h1798;
            14'd11111: out = 14'h1798;
            14'd11112: out = 14'h1797;
            14'd11113: out = 14'h1797;
            14'd11114: out = 14'h1796;
            14'd11115: out = 14'h1796;
            14'd11116: out = 14'h1795;
            14'd11117: out = 14'h1795;
            14'd11118: out = 14'h1794;
            14'd11119: out = 14'h1794;
            14'd11120: out = 14'h1793;
            14'd11121: out = 14'h1792;
            14'd11122: out = 14'h1792;
            14'd11123: out = 14'h1791;
            14'd11124: out = 14'h1791;
            14'd11125: out = 14'h1790;
            14'd11126: out = 14'h1790;
            14'd11127: out = 14'h178F;
            14'd11128: out = 14'h178F;
            14'd11129: out = 14'h178E;
            14'd11130: out = 14'h178E;
            14'd11131: out = 14'h178D;
            14'd11132: out = 14'h178C;
            14'd11133: out = 14'h178C;
            14'd11134: out = 14'h178B;
            14'd11135: out = 14'h178B;
            14'd11136: out = 14'h178A;
            14'd11137: out = 14'h178A;
            14'd11138: out = 14'h1789;
            14'd11139: out = 14'h1789;
            14'd11140: out = 14'h1788;
            14'd11141: out = 14'h1788;
            14'd11142: out = 14'h1787;
            14'd11143: out = 14'h1787;
            14'd11144: out = 14'h1786;
            14'd11145: out = 14'h1785;
            14'd11146: out = 14'h1785;
            14'd11147: out = 14'h1784;
            14'd11148: out = 14'h1784;
            14'd11149: out = 14'h1783;
            14'd11150: out = 14'h1783;
            14'd11151: out = 14'h1782;
            14'd11152: out = 14'h1782;
            14'd11153: out = 14'h1781;
            14'd11154: out = 14'h1781;
            14'd11155: out = 14'h1780;
            14'd11156: out = 14'h177F;
            14'd11157: out = 14'h177F;
            14'd11158: out = 14'h177E;
            14'd11159: out = 14'h177E;
            14'd11160: out = 14'h177D;
            14'd11161: out = 14'h177D;
            14'd11162: out = 14'h177C;
            14'd11163: out = 14'h177C;
            14'd11164: out = 14'h177B;
            14'd11165: out = 14'h177B;
            14'd11166: out = 14'h177A;
            14'd11167: out = 14'h177A;
            14'd11168: out = 14'h1779;
            14'd11169: out = 14'h1778;
            14'd11170: out = 14'h1778;
            14'd11171: out = 14'h1777;
            14'd11172: out = 14'h1777;
            14'd11173: out = 14'h1776;
            14'd11174: out = 14'h1776;
            14'd11175: out = 14'h1775;
            14'd11176: out = 14'h1775;
            14'd11177: out = 14'h1774;
            14'd11178: out = 14'h1774;
            14'd11179: out = 14'h1773;
            14'd11180: out = 14'h1773;
            14'd11181: out = 14'h1772;
            14'd11182: out = 14'h1772;
            14'd11183: out = 14'h1771;
            14'd11184: out = 14'h1770;
            14'd11185: out = 14'h1770;
            14'd11186: out = 14'h176F;
            14'd11187: out = 14'h176F;
            14'd11188: out = 14'h176E;
            14'd11189: out = 14'h176E;
            14'd11190: out = 14'h176D;
            14'd11191: out = 14'h176D;
            14'd11192: out = 14'h176C;
            14'd11193: out = 14'h176C;
            14'd11194: out = 14'h176B;
            14'd11195: out = 14'h176B;
            14'd11196: out = 14'h176A;
            14'd11197: out = 14'h1769;
            14'd11198: out = 14'h1769;
            14'd11199: out = 14'h1768;
            14'd11200: out = 14'h1768;
            14'd11201: out = 14'h1767;
            14'd11202: out = 14'h1767;
            14'd11203: out = 14'h1766;
            14'd11204: out = 14'h1766;
            14'd11205: out = 14'h1765;
            14'd11206: out = 14'h1765;
            14'd11207: out = 14'h1764;
            14'd11208: out = 14'h1764;
            14'd11209: out = 14'h1763;
            14'd11210: out = 14'h1763;
            14'd11211: out = 14'h1762;
            14'd11212: out = 14'h1761;
            14'd11213: out = 14'h1761;
            14'd11214: out = 14'h1760;
            14'd11215: out = 14'h1760;
            14'd11216: out = 14'h175F;
            14'd11217: out = 14'h175F;
            14'd11218: out = 14'h175E;
            14'd11219: out = 14'h175E;
            14'd11220: out = 14'h175D;
            14'd11221: out = 14'h175D;
            14'd11222: out = 14'h175C;
            14'd11223: out = 14'h175C;
            14'd11224: out = 14'h175B;
            14'd11225: out = 14'h175B;
            14'd11226: out = 14'h175A;
            14'd11227: out = 14'h1759;
            14'd11228: out = 14'h1759;
            14'd11229: out = 14'h1758;
            14'd11230: out = 14'h1758;
            14'd11231: out = 14'h1757;
            14'd11232: out = 14'h1757;
            14'd11233: out = 14'h1756;
            14'd11234: out = 14'h1756;
            14'd11235: out = 14'h1755;
            14'd11236: out = 14'h1755;
            14'd11237: out = 14'h1754;
            14'd11238: out = 14'h1754;
            14'd11239: out = 14'h1753;
            14'd11240: out = 14'h1753;
            14'd11241: out = 14'h1752;
            14'd11242: out = 14'h1751;
            14'd11243: out = 14'h1751;
            14'd11244: out = 14'h1750;
            14'd11245: out = 14'h1750;
            14'd11246: out = 14'h174F;
            14'd11247: out = 14'h174F;
            14'd11248: out = 14'h174E;
            14'd11249: out = 14'h174E;
            14'd11250: out = 14'h174D;
            14'd11251: out = 14'h174D;
            14'd11252: out = 14'h174C;
            14'd11253: out = 14'h174C;
            14'd11254: out = 14'h174B;
            14'd11255: out = 14'h174B;
            14'd11256: out = 14'h174A;
            14'd11257: out = 14'h174A;
            14'd11258: out = 14'h1749;
            14'd11259: out = 14'h1748;
            14'd11260: out = 14'h1748;
            14'd11261: out = 14'h1747;
            14'd11262: out = 14'h1747;
            14'd11263: out = 14'h1746;
            14'd11264: out = 14'h1746;
            14'd11265: out = 14'h1745;
            14'd11266: out = 14'h1745;
            14'd11267: out = 14'h1744;
            14'd11268: out = 14'h1744;
            14'd11269: out = 14'h1743;
            14'd11270: out = 14'h1743;
            14'd11271: out = 14'h1742;
            14'd11272: out = 14'h1742;
            14'd11273: out = 14'h1741;
            14'd11274: out = 14'h1741;
            14'd11275: out = 14'h1740;
            14'd11276: out = 14'h173F;
            14'd11277: out = 14'h173F;
            14'd11278: out = 14'h173E;
            14'd11279: out = 14'h173E;
            14'd11280: out = 14'h173D;
            14'd11281: out = 14'h173D;
            14'd11282: out = 14'h173C;
            14'd11283: out = 14'h173C;
            14'd11284: out = 14'h173B;
            14'd11285: out = 14'h173B;
            14'd11286: out = 14'h173A;
            14'd11287: out = 14'h173A;
            14'd11288: out = 14'h1739;
            14'd11289: out = 14'h1739;
            14'd11290: out = 14'h1738;
            14'd11291: out = 14'h1738;
            14'd11292: out = 14'h1737;
            14'd11293: out = 14'h1737;
            14'd11294: out = 14'h1736;
            14'd11295: out = 14'h1735;
            14'd11296: out = 14'h1735;
            14'd11297: out = 14'h1734;
            14'd11298: out = 14'h1734;
            14'd11299: out = 14'h1733;
            14'd11300: out = 14'h1733;
            14'd11301: out = 14'h1732;
            14'd11302: out = 14'h1732;
            14'd11303: out = 14'h1731;
            14'd11304: out = 14'h1731;
            14'd11305: out = 14'h1730;
            14'd11306: out = 14'h1730;
            14'd11307: out = 14'h172F;
            14'd11308: out = 14'h172F;
            14'd11309: out = 14'h172E;
            14'd11310: out = 14'h172E;
            14'd11311: out = 14'h172D;
            14'd11312: out = 14'h172D;
            14'd11313: out = 14'h172C;
            14'd11314: out = 14'h172B;
            14'd11315: out = 14'h172B;
            14'd11316: out = 14'h172A;
            14'd11317: out = 14'h172A;
            14'd11318: out = 14'h1729;
            14'd11319: out = 14'h1729;
            14'd11320: out = 14'h1728;
            14'd11321: out = 14'h1728;
            14'd11322: out = 14'h1727;
            14'd11323: out = 14'h1727;
            14'd11324: out = 14'h1726;
            14'd11325: out = 14'h1726;
            14'd11326: out = 14'h1725;
            14'd11327: out = 14'h1725;
            14'd11328: out = 14'h1724;
            14'd11329: out = 14'h1724;
            14'd11330: out = 14'h1723;
            14'd11331: out = 14'h1723;
            14'd11332: out = 14'h1722;
            14'd11333: out = 14'h1722;
            14'd11334: out = 14'h1721;
            14'd11335: out = 14'h1720;
            14'd11336: out = 14'h1720;
            14'd11337: out = 14'h171F;
            14'd11338: out = 14'h171F;
            14'd11339: out = 14'h171E;
            14'd11340: out = 14'h171E;
            14'd11341: out = 14'h171D;
            14'd11342: out = 14'h171D;
            14'd11343: out = 14'h171C;
            14'd11344: out = 14'h171C;
            14'd11345: out = 14'h171B;
            14'd11346: out = 14'h171B;
            14'd11347: out = 14'h171A;
            14'd11348: out = 14'h171A;
            14'd11349: out = 14'h1719;
            14'd11350: out = 14'h1719;
            14'd11351: out = 14'h1718;
            14'd11352: out = 14'h1718;
            14'd11353: out = 14'h1717;
            14'd11354: out = 14'h1717;
            14'd11355: out = 14'h1716;
            14'd11356: out = 14'h1716;
            14'd11357: out = 14'h1715;
            14'd11358: out = 14'h1715;
            14'd11359: out = 14'h1714;
            14'd11360: out = 14'h1713;
            14'd11361: out = 14'h1713;
            14'd11362: out = 14'h1712;
            14'd11363: out = 14'h1712;
            14'd11364: out = 14'h1711;
            14'd11365: out = 14'h1711;
            14'd11366: out = 14'h1710;
            14'd11367: out = 14'h1710;
            14'd11368: out = 14'h170F;
            14'd11369: out = 14'h170F;
            14'd11370: out = 14'h170E;
            14'd11371: out = 14'h170E;
            14'd11372: out = 14'h170D;
            14'd11373: out = 14'h170D;
            14'd11374: out = 14'h170C;
            14'd11375: out = 14'h170C;
            14'd11376: out = 14'h170B;
            14'd11377: out = 14'h170B;
            14'd11378: out = 14'h170A;
            14'd11379: out = 14'h170A;
            14'd11380: out = 14'h1709;
            14'd11381: out = 14'h1709;
            14'd11382: out = 14'h1708;
            14'd11383: out = 14'h1708;
            14'd11384: out = 14'h1707;
            14'd11385: out = 14'h1706;
            14'd11386: out = 14'h1706;
            14'd11387: out = 14'h1705;
            14'd11388: out = 14'h1705;
            14'd11389: out = 14'h1704;
            14'd11390: out = 14'h1704;
            14'd11391: out = 14'h1703;
            14'd11392: out = 14'h1703;
            14'd11393: out = 14'h1702;
            14'd11394: out = 14'h1702;
            14'd11395: out = 14'h1701;
            14'd11396: out = 14'h1701;
            14'd11397: out = 14'h1700;
            14'd11398: out = 14'h1700;
            14'd11399: out = 14'h16FF;
            14'd11400: out = 14'h16FF;
            14'd11401: out = 14'h16FE;
            14'd11402: out = 14'h16FE;
            14'd11403: out = 14'h16FD;
            14'd11404: out = 14'h16FD;
            14'd11405: out = 14'h16FC;
            14'd11406: out = 14'h16FC;
            14'd11407: out = 14'h16FB;
            14'd11408: out = 14'h16FB;
            14'd11409: out = 14'h16FA;
            14'd11410: out = 14'h16FA;
            14'd11411: out = 14'h16F9;
            14'd11412: out = 14'h16F9;
            14'd11413: out = 14'h16F8;
            14'd11414: out = 14'h16F8;
            14'd11415: out = 14'h16F7;
            14'd11416: out = 14'h16F6;
            14'd11417: out = 14'h16F6;
            14'd11418: out = 14'h16F5;
            14'd11419: out = 14'h16F5;
            14'd11420: out = 14'h16F4;
            14'd11421: out = 14'h16F4;
            14'd11422: out = 14'h16F3;
            14'd11423: out = 14'h16F3;
            14'd11424: out = 14'h16F2;
            14'd11425: out = 14'h16F2;
            14'd11426: out = 14'h16F1;
            14'd11427: out = 14'h16F1;
            14'd11428: out = 14'h16F0;
            14'd11429: out = 14'h16F0;
            14'd11430: out = 14'h16EF;
            14'd11431: out = 14'h16EF;
            14'd11432: out = 14'h16EE;
            14'd11433: out = 14'h16EE;
            14'd11434: out = 14'h16ED;
            14'd11435: out = 14'h16ED;
            14'd11436: out = 14'h16EC;
            14'd11437: out = 14'h16EC;
            14'd11438: out = 14'h16EB;
            14'd11439: out = 14'h16EB;
            14'd11440: out = 14'h16EA;
            14'd11441: out = 14'h16EA;
            14'd11442: out = 14'h16E9;
            14'd11443: out = 14'h16E9;
            14'd11444: out = 14'h16E8;
            14'd11445: out = 14'h16E8;
            14'd11446: out = 14'h16E7;
            14'd11447: out = 14'h16E7;
            14'd11448: out = 14'h16E6;
            14'd11449: out = 14'h16E6;
            14'd11450: out = 14'h16E5;
            14'd11451: out = 14'h16E5;
            14'd11452: out = 14'h16E4;
            14'd11453: out = 14'h16E4;
            14'd11454: out = 14'h16E3;
            14'd11455: out = 14'h16E2;
            14'd11456: out = 14'h16E2;
            14'd11457: out = 14'h16E1;
            14'd11458: out = 14'h16E1;
            14'd11459: out = 14'h16E0;
            14'd11460: out = 14'h16E0;
            14'd11461: out = 14'h16DF;
            14'd11462: out = 14'h16DF;
            14'd11463: out = 14'h16DE;
            14'd11464: out = 14'h16DE;
            14'd11465: out = 14'h16DD;
            14'd11466: out = 14'h16DD;
            14'd11467: out = 14'h16DC;
            14'd11468: out = 14'h16DC;
            14'd11469: out = 14'h16DB;
            14'd11470: out = 14'h16DB;
            14'd11471: out = 14'h16DA;
            14'd11472: out = 14'h16DA;
            14'd11473: out = 14'h16D9;
            14'd11474: out = 14'h16D9;
            14'd11475: out = 14'h16D8;
            14'd11476: out = 14'h16D8;
            14'd11477: out = 14'h16D7;
            14'd11478: out = 14'h16D7;
            14'd11479: out = 14'h16D6;
            14'd11480: out = 14'h16D6;
            14'd11481: out = 14'h16D5;
            14'd11482: out = 14'h16D5;
            14'd11483: out = 14'h16D4;
            14'd11484: out = 14'h16D4;
            14'd11485: out = 14'h16D3;
            14'd11486: out = 14'h16D3;
            14'd11487: out = 14'h16D2;
            14'd11488: out = 14'h16D2;
            14'd11489: out = 14'h16D1;
            14'd11490: out = 14'h16D1;
            14'd11491: out = 14'h16D0;
            14'd11492: out = 14'h16D0;
            14'd11493: out = 14'h16CF;
            14'd11494: out = 14'h16CF;
            14'd11495: out = 14'h16CE;
            14'd11496: out = 14'h16CE;
            14'd11497: out = 14'h16CD;
            14'd11498: out = 14'h16CD;
            14'd11499: out = 14'h16CC;
            14'd11500: out = 14'h16CC;
            14'd11501: out = 14'h16CB;
            14'd11502: out = 14'h16CB;
            14'd11503: out = 14'h16CA;
            14'd11504: out = 14'h16CA;
            14'd11505: out = 14'h16C9;
            14'd11506: out = 14'h16C9;
            14'd11507: out = 14'h16C8;
            14'd11508: out = 14'h16C7;
            14'd11509: out = 14'h16C7;
            14'd11510: out = 14'h16C6;
            14'd11511: out = 14'h16C6;
            14'd11512: out = 14'h16C5;
            14'd11513: out = 14'h16C5;
            14'd11514: out = 14'h16C4;
            14'd11515: out = 14'h16C4;
            14'd11516: out = 14'h16C3;
            14'd11517: out = 14'h16C3;
            14'd11518: out = 14'h16C2;
            14'd11519: out = 14'h16C2;
            14'd11520: out = 14'h16C1;
            14'd11521: out = 14'h16C1;
            14'd11522: out = 14'h16C0;
            14'd11523: out = 14'h16C0;
            14'd11524: out = 14'h16BF;
            14'd11525: out = 14'h16BF;
            14'd11526: out = 14'h16BE;
            14'd11527: out = 14'h16BE;
            14'd11528: out = 14'h16BD;
            14'd11529: out = 14'h16BD;
            14'd11530: out = 14'h16BC;
            14'd11531: out = 14'h16BC;
            14'd11532: out = 14'h16BB;
            14'd11533: out = 14'h16BB;
            14'd11534: out = 14'h16BA;
            14'd11535: out = 14'h16BA;
            14'd11536: out = 14'h16B9;
            14'd11537: out = 14'h16B9;
            14'd11538: out = 14'h16B8;
            14'd11539: out = 14'h16B8;
            14'd11540: out = 14'h16B7;
            14'd11541: out = 14'h16B7;
            14'd11542: out = 14'h16B6;
            14'd11543: out = 14'h16B6;
            14'd11544: out = 14'h16B5;
            14'd11545: out = 14'h16B5;
            14'd11546: out = 14'h16B4;
            14'd11547: out = 14'h16B4;
            14'd11548: out = 14'h16B3;
            14'd11549: out = 14'h16B3;
            14'd11550: out = 14'h16B2;
            14'd11551: out = 14'h16B2;
            14'd11552: out = 14'h16B1;
            14'd11553: out = 14'h16B1;
            14'd11554: out = 14'h16B0;
            14'd11555: out = 14'h16B0;
            14'd11556: out = 14'h16AF;
            14'd11557: out = 14'h16AF;
            14'd11558: out = 14'h16AE;
            14'd11559: out = 14'h16AE;
            14'd11560: out = 14'h16AD;
            14'd11561: out = 14'h16AD;
            14'd11562: out = 14'h16AC;
            14'd11563: out = 14'h16AC;
            14'd11564: out = 14'h16AB;
            14'd11565: out = 14'h16AB;
            14'd11566: out = 14'h16AA;
            14'd11567: out = 14'h16AA;
            14'd11568: out = 14'h16A9;
            14'd11569: out = 14'h16A9;
            14'd11570: out = 14'h16A8;
            14'd11571: out = 14'h16A8;
            14'd11572: out = 14'h16A7;
            14'd11573: out = 14'h16A7;
            14'd11574: out = 14'h16A6;
            14'd11575: out = 14'h16A6;
            14'd11576: out = 14'h16A5;
            14'd11577: out = 14'h16A5;
            14'd11578: out = 14'h16A4;
            14'd11579: out = 14'h16A4;
            14'd11580: out = 14'h16A3;
            14'd11581: out = 14'h16A3;
            14'd11582: out = 14'h16A2;
            14'd11583: out = 14'h16A2;
            14'd11584: out = 14'h16A1;
            14'd11585: out = 14'h16A1;
            14'd11586: out = 14'h16A0;
            14'd11587: out = 14'h16A0;
            14'd11588: out = 14'h169F;
            14'd11589: out = 14'h169F;
            14'd11590: out = 14'h169E;
            14'd11591: out = 14'h169E;
            14'd11592: out = 14'h169D;
            14'd11593: out = 14'h169D;
            14'd11594: out = 14'h169C;
            14'd11595: out = 14'h169C;
            14'd11596: out = 14'h169B;
            14'd11597: out = 14'h169B;
            14'd11598: out = 14'h169A;
            14'd11599: out = 14'h169A;
            14'd11600: out = 14'h1699;
            14'd11601: out = 14'h1699;
            14'd11602: out = 14'h1698;
            14'd11603: out = 14'h1698;
            14'd11604: out = 14'h1697;
            14'd11605: out = 14'h1697;
            14'd11606: out = 14'h1696;
            14'd11607: out = 14'h1696;
            14'd11608: out = 14'h1695;
            14'd11609: out = 14'h1695;
            14'd11610: out = 14'h1694;
            14'd11611: out = 14'h1694;
            14'd11612: out = 14'h1693;
            14'd11613: out = 14'h1693;
            14'd11614: out = 14'h1692;
            14'd11615: out = 14'h1692;
            14'd11616: out = 14'h1691;
            14'd11617: out = 14'h1691;
            14'd11618: out = 14'h1690;
            14'd11619: out = 14'h1690;
            14'd11620: out = 14'h168F;
            14'd11621: out = 14'h168F;
            14'd11622: out = 14'h168E;
            14'd11623: out = 14'h168E;
            14'd11624: out = 14'h168D;
            14'd11625: out = 14'h168D;
            14'd11626: out = 14'h168C;
            14'd11627: out = 14'h168C;
            14'd11628: out = 14'h168B;
            14'd11629: out = 14'h168B;
            14'd11630: out = 14'h168A;
            14'd11631: out = 14'h168A;
            14'd11632: out = 14'h1689;
            14'd11633: out = 14'h1689;
            14'd11634: out = 14'h1688;
            14'd11635: out = 14'h1688;
            14'd11636: out = 14'h1687;
            14'd11637: out = 14'h1687;
            14'd11638: out = 14'h1686;
            14'd11639: out = 14'h1686;
            14'd11640: out = 14'h1685;
            14'd11641: out = 14'h1685;
            14'd11642: out = 14'h1684;
            14'd11643: out = 14'h1684;
            14'd11644: out = 14'h1683;
            14'd11645: out = 14'h1683;
            14'd11646: out = 14'h1682;
            14'd11647: out = 14'h1682;
            14'd11648: out = 14'h1681;
            14'd11649: out = 14'h1681;
            14'd11650: out = 14'h1680;
            14'd11651: out = 14'h1680;
            14'd11652: out = 14'h167F;
            14'd11653: out = 14'h167F;
            14'd11654: out = 14'h167E;
            14'd11655: out = 14'h167E;
            14'd11656: out = 14'h167D;
            14'd11657: out = 14'h167D;
            14'd11658: out = 14'h167C;
            14'd11659: out = 14'h167C;
            14'd11660: out = 14'h167B;
            14'd11661: out = 14'h167B;
            14'd11662: out = 14'h167A;
            14'd11663: out = 14'h167A;
            14'd11664: out = 14'h167A;
            14'd11665: out = 14'h1679;
            14'd11666: out = 14'h1679;
            14'd11667: out = 14'h1678;
            14'd11668: out = 14'h1678;
            14'd11669: out = 14'h1677;
            14'd11670: out = 14'h1677;
            14'd11671: out = 14'h1676;
            14'd11672: out = 14'h1676;
            14'd11673: out = 14'h1675;
            14'd11674: out = 14'h1675;
            14'd11675: out = 14'h1674;
            14'd11676: out = 14'h1674;
            14'd11677: out = 14'h1673;
            14'd11678: out = 14'h1673;
            14'd11679: out = 14'h1672;
            14'd11680: out = 14'h1672;
            14'd11681: out = 14'h1671;
            14'd11682: out = 14'h1671;
            14'd11683: out = 14'h1670;
            14'd11684: out = 14'h1670;
            14'd11685: out = 14'h166F;
            14'd11686: out = 14'h166F;
            14'd11687: out = 14'h166E;
            14'd11688: out = 14'h166E;
            14'd11689: out = 14'h166D;
            14'd11690: out = 14'h166D;
            14'd11691: out = 14'h166C;
            14'd11692: out = 14'h166C;
            14'd11693: out = 14'h166B;
            14'd11694: out = 14'h166B;
            14'd11695: out = 14'h166A;
            14'd11696: out = 14'h166A;
            14'd11697: out = 14'h1669;
            14'd11698: out = 14'h1669;
            14'd11699: out = 14'h1668;
            14'd11700: out = 14'h1668;
            14'd11701: out = 14'h1667;
            14'd11702: out = 14'h1667;
            14'd11703: out = 14'h1666;
            14'd11704: out = 14'h1666;
            14'd11705: out = 14'h1665;
            14'd11706: out = 14'h1665;
            14'd11707: out = 14'h1664;
            14'd11708: out = 14'h1664;
            14'd11709: out = 14'h1663;
            14'd11710: out = 14'h1663;
            14'd11711: out = 14'h1662;
            14'd11712: out = 14'h1662;
            14'd11713: out = 14'h1661;
            14'd11714: out = 14'h1661;
            14'd11715: out = 14'h1660;
            14'd11716: out = 14'h1660;
            14'd11717: out = 14'h165F;
            14'd11718: out = 14'h165F;
            14'd11719: out = 14'h165F;
            14'd11720: out = 14'h165E;
            14'd11721: out = 14'h165E;
            14'd11722: out = 14'h165D;
            14'd11723: out = 14'h165D;
            14'd11724: out = 14'h165C;
            14'd11725: out = 14'h165C;
            14'd11726: out = 14'h165B;
            14'd11727: out = 14'h165B;
            14'd11728: out = 14'h165A;
            14'd11729: out = 14'h165A;
            14'd11730: out = 14'h1659;
            14'd11731: out = 14'h1659;
            14'd11732: out = 14'h1658;
            14'd11733: out = 14'h1658;
            14'd11734: out = 14'h1657;
            14'd11735: out = 14'h1657;
            14'd11736: out = 14'h1656;
            14'd11737: out = 14'h1656;
            14'd11738: out = 14'h1655;
            14'd11739: out = 14'h1655;
            14'd11740: out = 14'h1654;
            14'd11741: out = 14'h1654;
            14'd11742: out = 14'h1653;
            14'd11743: out = 14'h1653;
            14'd11744: out = 14'h1652;
            14'd11745: out = 14'h1652;
            14'd11746: out = 14'h1651;
            14'd11747: out = 14'h1651;
            14'd11748: out = 14'h1650;
            14'd11749: out = 14'h1650;
            14'd11750: out = 14'h164F;
            14'd11751: out = 14'h164F;
            14'd11752: out = 14'h164E;
            14'd11753: out = 14'h164E;
            14'd11754: out = 14'h164D;
            14'd11755: out = 14'h164D;
            14'd11756: out = 14'h164C;
            14'd11757: out = 14'h164C;
            14'd11758: out = 14'h164C;
            14'd11759: out = 14'h164B;
            14'd11760: out = 14'h164B;
            14'd11761: out = 14'h164A;
            14'd11762: out = 14'h164A;
            14'd11763: out = 14'h1649;
            14'd11764: out = 14'h1649;
            14'd11765: out = 14'h1648;
            14'd11766: out = 14'h1648;
            14'd11767: out = 14'h1647;
            14'd11768: out = 14'h1647;
            14'd11769: out = 14'h1646;
            14'd11770: out = 14'h1646;
            14'd11771: out = 14'h1645;
            14'd11772: out = 14'h1645;
            14'd11773: out = 14'h1644;
            14'd11774: out = 14'h1644;
            14'd11775: out = 14'h1643;
            14'd11776: out = 14'h1643;
            14'd11777: out = 14'h1642;
            14'd11778: out = 14'h1642;
            14'd11779: out = 14'h1641;
            14'd11780: out = 14'h1641;
            14'd11781: out = 14'h1640;
            14'd11782: out = 14'h1640;
            14'd11783: out = 14'h163F;
            14'd11784: out = 14'h163F;
            14'd11785: out = 14'h163E;
            14'd11786: out = 14'h163E;
            14'd11787: out = 14'h163D;
            14'd11788: out = 14'h163D;
            14'd11789: out = 14'h163C;
            14'd11790: out = 14'h163C;
            14'd11791: out = 14'h163C;
            14'd11792: out = 14'h163B;
            14'd11793: out = 14'h163B;
            14'd11794: out = 14'h163A;
            14'd11795: out = 14'h163A;
            14'd11796: out = 14'h1639;
            14'd11797: out = 14'h1639;
            14'd11798: out = 14'h1638;
            14'd11799: out = 14'h1638;
            14'd11800: out = 14'h1637;
            14'd11801: out = 14'h1637;
            14'd11802: out = 14'h1636;
            14'd11803: out = 14'h1636;
            14'd11804: out = 14'h1635;
            14'd11805: out = 14'h1635;
            14'd11806: out = 14'h1634;
            14'd11807: out = 14'h1634;
            14'd11808: out = 14'h1633;
            14'd11809: out = 14'h1633;
            14'd11810: out = 14'h1632;
            14'd11811: out = 14'h1632;
            14'd11812: out = 14'h1631;
            14'd11813: out = 14'h1631;
            14'd11814: out = 14'h1630;
            14'd11815: out = 14'h1630;
            14'd11816: out = 14'h162F;
            14'd11817: out = 14'h162F;
            14'd11818: out = 14'h162F;
            14'd11819: out = 14'h162E;
            14'd11820: out = 14'h162E;
            14'd11821: out = 14'h162D;
            14'd11822: out = 14'h162D;
            14'd11823: out = 14'h162C;
            14'd11824: out = 14'h162C;
            14'd11825: out = 14'h162B;
            14'd11826: out = 14'h162B;
            14'd11827: out = 14'h162A;
            14'd11828: out = 14'h162A;
            14'd11829: out = 14'h1629;
            14'd11830: out = 14'h1629;
            14'd11831: out = 14'h1628;
            14'd11832: out = 14'h1628;
            14'd11833: out = 14'h1627;
            14'd11834: out = 14'h1627;
            14'd11835: out = 14'h1626;
            14'd11836: out = 14'h1626;
            14'd11837: out = 14'h1625;
            14'd11838: out = 14'h1625;
            14'd11839: out = 14'h1624;
            14'd11840: out = 14'h1624;
            14'd11841: out = 14'h1623;
            14'd11842: out = 14'h1623;
            14'd11843: out = 14'h1623;
            14'd11844: out = 14'h1622;
            14'd11845: out = 14'h1622;
            14'd11846: out = 14'h1621;
            14'd11847: out = 14'h1621;
            14'd11848: out = 14'h1620;
            14'd11849: out = 14'h1620;
            14'd11850: out = 14'h161F;
            14'd11851: out = 14'h161F;
            14'd11852: out = 14'h161E;
            14'd11853: out = 14'h161E;
            14'd11854: out = 14'h161D;
            14'd11855: out = 14'h161D;
            14'd11856: out = 14'h161C;
            14'd11857: out = 14'h161C;
            14'd11858: out = 14'h161B;
            14'd11859: out = 14'h161B;
            14'd11860: out = 14'h161A;
            14'd11861: out = 14'h161A;
            14'd11862: out = 14'h1619;
            14'd11863: out = 14'h1619;
            14'd11864: out = 14'h1619;
            14'd11865: out = 14'h1618;
            14'd11866: out = 14'h1618;
            14'd11867: out = 14'h1617;
            14'd11868: out = 14'h1617;
            14'd11869: out = 14'h1616;
            14'd11870: out = 14'h1616;
            14'd11871: out = 14'h1615;
            14'd11872: out = 14'h1615;
            14'd11873: out = 14'h1614;
            14'd11874: out = 14'h1614;
            14'd11875: out = 14'h1613;
            14'd11876: out = 14'h1613;
            14'd11877: out = 14'h1612;
            14'd11878: out = 14'h1612;
            14'd11879: out = 14'h1611;
            14'd11880: out = 14'h1611;
            14'd11881: out = 14'h1610;
            14'd11882: out = 14'h1610;
            14'd11883: out = 14'h160F;
            14'd11884: out = 14'h160F;
            14'd11885: out = 14'h160F;
            14'd11886: out = 14'h160E;
            14'd11887: out = 14'h160E;
            14'd11888: out = 14'h160D;
            14'd11889: out = 14'h160D;
            14'd11890: out = 14'h160C;
            14'd11891: out = 14'h160C;
            14'd11892: out = 14'h160B;
            14'd11893: out = 14'h160B;
            14'd11894: out = 14'h160A;
            14'd11895: out = 14'h160A;
            14'd11896: out = 14'h1609;
            14'd11897: out = 14'h1609;
            14'd11898: out = 14'h1608;
            14'd11899: out = 14'h1608;
            14'd11900: out = 14'h1607;
            14'd11901: out = 14'h1607;
            14'd11902: out = 14'h1606;
            14'd11903: out = 14'h1606;
            14'd11904: out = 14'h1606;
            14'd11905: out = 14'h1605;
            14'd11906: out = 14'h1605;
            14'd11907: out = 14'h1604;
            14'd11908: out = 14'h1604;
            14'd11909: out = 14'h1603;
            14'd11910: out = 14'h1603;
            14'd11911: out = 14'h1602;
            14'd11912: out = 14'h1602;
            14'd11913: out = 14'h1601;
            14'd11914: out = 14'h1601;
            14'd11915: out = 14'h1600;
            14'd11916: out = 14'h1600;
            14'd11917: out = 14'h15FF;
            14'd11918: out = 14'h15FF;
            14'd11919: out = 14'h15FE;
            14'd11920: out = 14'h15FE;
            14'd11921: out = 14'h15FD;
            14'd11922: out = 14'h15FD;
            14'd11923: out = 14'h15FD;
            14'd11924: out = 14'h15FC;
            14'd11925: out = 14'h15FC;
            14'd11926: out = 14'h15FB;
            14'd11927: out = 14'h15FB;
            14'd11928: out = 14'h15FA;
            14'd11929: out = 14'h15FA;
            14'd11930: out = 14'h15F9;
            14'd11931: out = 14'h15F9;
            14'd11932: out = 14'h15F8;
            14'd11933: out = 14'h15F8;
            14'd11934: out = 14'h15F7;
            14'd11935: out = 14'h15F7;
            14'd11936: out = 14'h15F6;
            14'd11937: out = 14'h15F6;
            14'd11938: out = 14'h15F5;
            14'd11939: out = 14'h15F5;
            14'd11940: out = 14'h15F5;
            14'd11941: out = 14'h15F4;
            14'd11942: out = 14'h15F4;
            14'd11943: out = 14'h15F3;
            14'd11944: out = 14'h15F3;
            14'd11945: out = 14'h15F2;
            14'd11946: out = 14'h15F2;
            14'd11947: out = 14'h15F1;
            14'd11948: out = 14'h15F1;
            14'd11949: out = 14'h15F0;
            14'd11950: out = 14'h15F0;
            14'd11951: out = 14'h15EF;
            14'd11952: out = 14'h15EF;
            14'd11953: out = 14'h15EE;
            14'd11954: out = 14'h15EE;
            14'd11955: out = 14'h15ED;
            14'd11956: out = 14'h15ED;
            14'd11957: out = 14'h15ED;
            14'd11958: out = 14'h15EC;
            14'd11959: out = 14'h15EC;
            14'd11960: out = 14'h15EB;
            14'd11961: out = 14'h15EB;
            14'd11962: out = 14'h15EA;
            14'd11963: out = 14'h15EA;
            14'd11964: out = 14'h15E9;
            14'd11965: out = 14'h15E9;
            14'd11966: out = 14'h15E8;
            14'd11967: out = 14'h15E8;
            14'd11968: out = 14'h15E7;
            14'd11969: out = 14'h15E7;
            14'd11970: out = 14'h15E6;
            14'd11971: out = 14'h15E6;
            14'd11972: out = 14'h15E5;
            14'd11973: out = 14'h15E5;
            14'd11974: out = 14'h15E5;
            14'd11975: out = 14'h15E4;
            14'd11976: out = 14'h15E4;
            14'd11977: out = 14'h15E3;
            14'd11978: out = 14'h15E3;
            14'd11979: out = 14'h15E2;
            14'd11980: out = 14'h15E2;
            14'd11981: out = 14'h15E1;
            14'd11982: out = 14'h15E1;
            14'd11983: out = 14'h15E0;
            14'd11984: out = 14'h15E0;
            14'd11985: out = 14'h15DF;
            14'd11986: out = 14'h15DF;
            14'd11987: out = 14'h15DE;
            14'd11988: out = 14'h15DE;
            14'd11989: out = 14'h15DE;
            14'd11990: out = 14'h15DD;
            14'd11991: out = 14'h15DD;
            14'd11992: out = 14'h15DC;
            14'd11993: out = 14'h15DC;
            14'd11994: out = 14'h15DB;
            14'd11995: out = 14'h15DB;
            14'd11996: out = 14'h15DA;
            14'd11997: out = 14'h15DA;
            14'd11998: out = 14'h15D9;
            14'd11999: out = 14'h15D9;
            14'd12000: out = 14'h15D8;
            14'd12001: out = 14'h15D8;
            14'd12002: out = 14'h15D7;
            14'd12003: out = 14'h15D7;
            14'd12004: out = 14'h15D7;
            14'd12005: out = 14'h15D6;
            14'd12006: out = 14'h15D6;
            14'd12007: out = 14'h15D5;
            14'd12008: out = 14'h15D5;
            14'd12009: out = 14'h15D4;
            14'd12010: out = 14'h15D4;
            14'd12011: out = 14'h15D3;
            14'd12012: out = 14'h15D3;
            14'd12013: out = 14'h15D2;
            14'd12014: out = 14'h15D2;
            14'd12015: out = 14'h15D1;
            14'd12016: out = 14'h15D1;
            14'd12017: out = 14'h15D0;
            14'd12018: out = 14'h15D0;
            14'd12019: out = 14'h15D0;
            14'd12020: out = 14'h15CF;
            14'd12021: out = 14'h15CF;
            14'd12022: out = 14'h15CE;
            14'd12023: out = 14'h15CE;
            14'd12024: out = 14'h15CD;
            14'd12025: out = 14'h15CD;
            14'd12026: out = 14'h15CC;
            14'd12027: out = 14'h15CC;
            14'd12028: out = 14'h15CB;
            14'd12029: out = 14'h15CB;
            14'd12030: out = 14'h15CA;
            14'd12031: out = 14'h15CA;
            14'd12032: out = 14'h15CA;
            14'd12033: out = 14'h15C9;
            14'd12034: out = 14'h15C9;
            14'd12035: out = 14'h15C8;
            14'd12036: out = 14'h15C8;
            14'd12037: out = 14'h15C7;
            14'd12038: out = 14'h15C7;
            14'd12039: out = 14'h15C6;
            14'd12040: out = 14'h15C6;
            14'd12041: out = 14'h15C5;
            14'd12042: out = 14'h15C5;
            14'd12043: out = 14'h15C4;
            14'd12044: out = 14'h15C4;
            14'd12045: out = 14'h15C4;
            14'd12046: out = 14'h15C3;
            14'd12047: out = 14'h15C3;
            14'd12048: out = 14'h15C2;
            14'd12049: out = 14'h15C2;
            14'd12050: out = 14'h15C1;
            14'd12051: out = 14'h15C1;
            14'd12052: out = 14'h15C0;
            14'd12053: out = 14'h15C0;
            14'd12054: out = 14'h15BF;
            14'd12055: out = 14'h15BF;
            14'd12056: out = 14'h15BE;
            14'd12057: out = 14'h15BE;
            14'd12058: out = 14'h15BE;
            14'd12059: out = 14'h15BD;
            14'd12060: out = 14'h15BD;
            14'd12061: out = 14'h15BC;
            14'd12062: out = 14'h15BC;
            14'd12063: out = 14'h15BB;
            14'd12064: out = 14'h15BB;
            14'd12065: out = 14'h15BA;
            14'd12066: out = 14'h15BA;
            14'd12067: out = 14'h15B9;
            14'd12068: out = 14'h15B9;
            14'd12069: out = 14'h15B8;
            14'd12070: out = 14'h15B8;
            14'd12071: out = 14'h15B8;
            14'd12072: out = 14'h15B7;
            14'd12073: out = 14'h15B7;
            14'd12074: out = 14'h15B6;
            14'd12075: out = 14'h15B6;
            14'd12076: out = 14'h15B5;
            14'd12077: out = 14'h15B5;
            14'd12078: out = 14'h15B4;
            14'd12079: out = 14'h15B4;
            14'd12080: out = 14'h15B3;
            14'd12081: out = 14'h15B3;
            14'd12082: out = 14'h15B2;
            14'd12083: out = 14'h15B2;
            14'd12084: out = 14'h15B2;
            14'd12085: out = 14'h15B1;
            14'd12086: out = 14'h15B1;
            14'd12087: out = 14'h15B0;
            14'd12088: out = 14'h15B0;
            14'd12089: out = 14'h15AF;
            14'd12090: out = 14'h15AF;
            14'd12091: out = 14'h15AE;
            14'd12092: out = 14'h15AE;
            14'd12093: out = 14'h15AD;
            14'd12094: out = 14'h15AD;
            14'd12095: out = 14'h15AC;
            14'd12096: out = 14'h15AC;
            14'd12097: out = 14'h15AC;
            14'd12098: out = 14'h15AB;
            14'd12099: out = 14'h15AB;
            14'd12100: out = 14'h15AA;
            14'd12101: out = 14'h15AA;
            14'd12102: out = 14'h15A9;
            14'd12103: out = 14'h15A9;
            14'd12104: out = 14'h15A8;
            14'd12105: out = 14'h15A8;
            14'd12106: out = 14'h15A7;
            14'd12107: out = 14'h15A7;
            14'd12108: out = 14'h15A7;
            14'd12109: out = 14'h15A6;
            14'd12110: out = 14'h15A6;
            14'd12111: out = 14'h15A5;
            14'd12112: out = 14'h15A5;
            14'd12113: out = 14'h15A4;
            14'd12114: out = 14'h15A4;
            14'd12115: out = 14'h15A3;
            14'd12116: out = 14'h15A3;
            14'd12117: out = 14'h15A2;
            14'd12118: out = 14'h15A2;
            14'd12119: out = 14'h15A1;
            14'd12120: out = 14'h15A1;
            14'd12121: out = 14'h15A1;
            14'd12122: out = 14'h15A0;
            14'd12123: out = 14'h15A0;
            14'd12124: out = 14'h159F;
            14'd12125: out = 14'h159F;
            14'd12126: out = 14'h159E;
            14'd12127: out = 14'h159E;
            14'd12128: out = 14'h159D;
            14'd12129: out = 14'h159D;
            14'd12130: out = 14'h159C;
            14'd12131: out = 14'h159C;
            14'd12132: out = 14'h159C;
            14'd12133: out = 14'h159B;
            14'd12134: out = 14'h159B;
            14'd12135: out = 14'h159A;
            14'd12136: out = 14'h159A;
            14'd12137: out = 14'h1599;
            14'd12138: out = 14'h1599;
            14'd12139: out = 14'h1598;
            14'd12140: out = 14'h1598;
            14'd12141: out = 14'h1597;
            14'd12142: out = 14'h1597;
            14'd12143: out = 14'h1597;
            14'd12144: out = 14'h1596;
            14'd12145: out = 14'h1596;
            14'd12146: out = 14'h1595;
            14'd12147: out = 14'h1595;
            14'd12148: out = 14'h1594;
            14'd12149: out = 14'h1594;
            14'd12150: out = 14'h1593;
            14'd12151: out = 14'h1593;
            14'd12152: out = 14'h1592;
            14'd12153: out = 14'h1592;
            14'd12154: out = 14'h1592;
            14'd12155: out = 14'h1591;
            14'd12156: out = 14'h1591;
            14'd12157: out = 14'h1590;
            14'd12158: out = 14'h1590;
            14'd12159: out = 14'h158F;
            14'd12160: out = 14'h158F;
            14'd12161: out = 14'h158E;
            14'd12162: out = 14'h158E;
            14'd12163: out = 14'h158D;
            14'd12164: out = 14'h158D;
            14'd12165: out = 14'h158D;
            14'd12166: out = 14'h158C;
            14'd12167: out = 14'h158C;
            14'd12168: out = 14'h158B;
            14'd12169: out = 14'h158B;
            14'd12170: out = 14'h158A;
            14'd12171: out = 14'h158A;
            14'd12172: out = 14'h1589;
            14'd12173: out = 14'h1589;
            14'd12174: out = 14'h1588;
            14'd12175: out = 14'h1588;
            14'd12176: out = 14'h1588;
            14'd12177: out = 14'h1587;
            14'd12178: out = 14'h1587;
            14'd12179: out = 14'h1586;
            14'd12180: out = 14'h1586;
            14'd12181: out = 14'h1585;
            14'd12182: out = 14'h1585;
            14'd12183: out = 14'h1584;
            14'd12184: out = 14'h1584;
            14'd12185: out = 14'h1583;
            14'd12186: out = 14'h1583;
            14'd12187: out = 14'h1583;
            14'd12188: out = 14'h1582;
            14'd12189: out = 14'h1582;
            14'd12190: out = 14'h1581;
            14'd12191: out = 14'h1581;
            14'd12192: out = 14'h1580;
            14'd12193: out = 14'h1580;
            14'd12194: out = 14'h157F;
            14'd12195: out = 14'h157F;
            14'd12196: out = 14'h157F;
            14'd12197: out = 14'h157E;
            14'd12198: out = 14'h157E;
            14'd12199: out = 14'h157D;
            14'd12200: out = 14'h157D;
            14'd12201: out = 14'h157C;
            14'd12202: out = 14'h157C;
            14'd12203: out = 14'h157B;
            14'd12204: out = 14'h157B;
            14'd12205: out = 14'h157A;
            14'd12206: out = 14'h157A;
            14'd12207: out = 14'h157A;
            14'd12208: out = 14'h1579;
            14'd12209: out = 14'h1579;
            14'd12210: out = 14'h1578;
            14'd12211: out = 14'h1578;
            14'd12212: out = 14'h1577;
            14'd12213: out = 14'h1577;
            14'd12214: out = 14'h1576;
            14'd12215: out = 14'h1576;
            14'd12216: out = 14'h1576;
            14'd12217: out = 14'h1575;
            14'd12218: out = 14'h1575;
            14'd12219: out = 14'h1574;
            14'd12220: out = 14'h1574;
            14'd12221: out = 14'h1573;
            14'd12222: out = 14'h1573;
            14'd12223: out = 14'h1572;
            14'd12224: out = 14'h1572;
            14'd12225: out = 14'h1571;
            14'd12226: out = 14'h1571;
            14'd12227: out = 14'h1571;
            14'd12228: out = 14'h1570;
            14'd12229: out = 14'h1570;
            14'd12230: out = 14'h156F;
            14'd12231: out = 14'h156F;
            14'd12232: out = 14'h156E;
            14'd12233: out = 14'h156E;
            14'd12234: out = 14'h156D;
            14'd12235: out = 14'h156D;
            14'd12236: out = 14'h156D;
            14'd12237: out = 14'h156C;
            14'd12238: out = 14'h156C;
            14'd12239: out = 14'h156B;
            14'd12240: out = 14'h156B;
            14'd12241: out = 14'h156A;
            14'd12242: out = 14'h156A;
            14'd12243: out = 14'h1569;
            14'd12244: out = 14'h1569;
            14'd12245: out = 14'h1569;
            14'd12246: out = 14'h1568;
            14'd12247: out = 14'h1568;
            14'd12248: out = 14'h1567;
            14'd12249: out = 14'h1567;
            14'd12250: out = 14'h1566;
            14'd12251: out = 14'h1566;
            14'd12252: out = 14'h1565;
            14'd12253: out = 14'h1565;
            14'd12254: out = 14'h1564;
            14'd12255: out = 14'h1564;
            14'd12256: out = 14'h1564;
            14'd12257: out = 14'h1563;
            14'd12258: out = 14'h1563;
            14'd12259: out = 14'h1562;
            14'd12260: out = 14'h1562;
            14'd12261: out = 14'h1561;
            14'd12262: out = 14'h1561;
            14'd12263: out = 14'h1560;
            14'd12264: out = 14'h1560;
            14'd12265: out = 14'h1560;
            14'd12266: out = 14'h155F;
            14'd12267: out = 14'h155F;
            14'd12268: out = 14'h155E;
            14'd12269: out = 14'h155E;
            14'd12270: out = 14'h155D;
            14'd12271: out = 14'h155D;
            14'd12272: out = 14'h155C;
            14'd12273: out = 14'h155C;
            14'd12274: out = 14'h155C;
            14'd12275: out = 14'h155B;
            14'd12276: out = 14'h155B;
            14'd12277: out = 14'h155A;
            14'd12278: out = 14'h155A;
            14'd12279: out = 14'h1559;
            14'd12280: out = 14'h1559;
            14'd12281: out = 14'h1558;
            14'd12282: out = 14'h1558;
            14'd12283: out = 14'h1558;
            14'd12284: out = 14'h1557;
            14'd12285: out = 14'h1557;
            14'd12286: out = 14'h1556;
            14'd12287: out = 14'h1556;
            14'd12288: out = 14'h1555;
            14'd12289: out = 14'h1555;
            14'd12290: out = 14'h1554;
            14'd12291: out = 14'h1554;
            14'd12292: out = 14'h1554;
            14'd12293: out = 14'h1553;
            14'd12294: out = 14'h1553;
            14'd12295: out = 14'h1552;
            14'd12296: out = 14'h1552;
            14'd12297: out = 14'h1551;
            14'd12298: out = 14'h1551;
            14'd12299: out = 14'h1550;
            14'd12300: out = 14'h1550;
            14'd12301: out = 14'h1550;
            14'd12302: out = 14'h154F;
            14'd12303: out = 14'h154F;
            14'd12304: out = 14'h154E;
            14'd12305: out = 14'h154E;
            14'd12306: out = 14'h154D;
            14'd12307: out = 14'h154D;
            14'd12308: out = 14'h154C;
            14'd12309: out = 14'h154C;
            14'd12310: out = 14'h154C;
            14'd12311: out = 14'h154B;
            14'd12312: out = 14'h154B;
            14'd12313: out = 14'h154A;
            14'd12314: out = 14'h154A;
            14'd12315: out = 14'h1549;
            14'd12316: out = 14'h1549;
            14'd12317: out = 14'h1548;
            14'd12318: out = 14'h1548;
            14'd12319: out = 14'h1548;
            14'd12320: out = 14'h1547;
            14'd12321: out = 14'h1547;
            14'd12322: out = 14'h1546;
            14'd12323: out = 14'h1546;
            14'd12324: out = 14'h1545;
            14'd12325: out = 14'h1545;
            14'd12326: out = 14'h1544;
            14'd12327: out = 14'h1544;
            14'd12328: out = 14'h1544;
            14'd12329: out = 14'h1543;
            14'd12330: out = 14'h1543;
            14'd12331: out = 14'h1542;
            14'd12332: out = 14'h1542;
            14'd12333: out = 14'h1541;
            14'd12334: out = 14'h1541;
            14'd12335: out = 14'h1541;
            14'd12336: out = 14'h1540;
            14'd12337: out = 14'h1540;
            14'd12338: out = 14'h153F;
            14'd12339: out = 14'h153F;
            14'd12340: out = 14'h153E;
            14'd12341: out = 14'h153E;
            14'd12342: out = 14'h153D;
            14'd12343: out = 14'h153D;
            14'd12344: out = 14'h153D;
            14'd12345: out = 14'h153C;
            14'd12346: out = 14'h153C;
            14'd12347: out = 14'h153B;
            14'd12348: out = 14'h153B;
            14'd12349: out = 14'h153A;
            14'd12350: out = 14'h153A;
            14'd12351: out = 14'h1539;
            14'd12352: out = 14'h1539;
            14'd12353: out = 14'h1539;
            14'd12354: out = 14'h1538;
            14'd12355: out = 14'h1538;
            14'd12356: out = 14'h1537;
            14'd12357: out = 14'h1537;
            14'd12358: out = 14'h1536;
            14'd12359: out = 14'h1536;
            14'd12360: out = 14'h1536;
            14'd12361: out = 14'h1535;
            14'd12362: out = 14'h1535;
            14'd12363: out = 14'h1534;
            14'd12364: out = 14'h1534;
            14'd12365: out = 14'h1533;
            14'd12366: out = 14'h1533;
            14'd12367: out = 14'h1532;
            14'd12368: out = 14'h1532;
            14'd12369: out = 14'h1532;
            14'd12370: out = 14'h1531;
            14'd12371: out = 14'h1531;
            14'd12372: out = 14'h1530;
            14'd12373: out = 14'h1530;
            14'd12374: out = 14'h152F;
            14'd12375: out = 14'h152F;
            14'd12376: out = 14'h152F;
            14'd12377: out = 14'h152E;
            14'd12378: out = 14'h152E;
            14'd12379: out = 14'h152D;
            14'd12380: out = 14'h152D;
            14'd12381: out = 14'h152C;
            14'd12382: out = 14'h152C;
            14'd12383: out = 14'h152B;
            14'd12384: out = 14'h152B;
            14'd12385: out = 14'h152B;
            14'd12386: out = 14'h152A;
            14'd12387: out = 14'h152A;
            14'd12388: out = 14'h1529;
            14'd12389: out = 14'h1529;
            14'd12390: out = 14'h1528;
            14'd12391: out = 14'h1528;
            14'd12392: out = 14'h1527;
            14'd12393: out = 14'h1527;
            14'd12394: out = 14'h1527;
            14'd12395: out = 14'h1526;
            14'd12396: out = 14'h1526;
            14'd12397: out = 14'h1525;
            14'd12398: out = 14'h1525;
            14'd12399: out = 14'h1524;
            14'd12400: out = 14'h1524;
            14'd12401: out = 14'h1524;
            14'd12402: out = 14'h1523;
            14'd12403: out = 14'h1523;
            14'd12404: out = 14'h1522;
            14'd12405: out = 14'h1522;
            14'd12406: out = 14'h1521;
            14'd12407: out = 14'h1521;
            14'd12408: out = 14'h1521;
            14'd12409: out = 14'h1520;
            14'd12410: out = 14'h1520;
            14'd12411: out = 14'h151F;
            14'd12412: out = 14'h151F;
            14'd12413: out = 14'h151E;
            14'd12414: out = 14'h151E;
            14'd12415: out = 14'h151D;
            14'd12416: out = 14'h151D;
            14'd12417: out = 14'h151D;
            14'd12418: out = 14'h151C;
            14'd12419: out = 14'h151C;
            14'd12420: out = 14'h151B;
            14'd12421: out = 14'h151B;
            14'd12422: out = 14'h151A;
            14'd12423: out = 14'h151A;
            14'd12424: out = 14'h151A;
            14'd12425: out = 14'h1519;
            14'd12426: out = 14'h1519;
            14'd12427: out = 14'h1518;
            14'd12428: out = 14'h1518;
            14'd12429: out = 14'h1517;
            14'd12430: out = 14'h1517;
            14'd12431: out = 14'h1517;
            14'd12432: out = 14'h1516;
            14'd12433: out = 14'h1516;
            14'd12434: out = 14'h1515;
            14'd12435: out = 14'h1515;
            14'd12436: out = 14'h1514;
            14'd12437: out = 14'h1514;
            14'd12438: out = 14'h1513;
            14'd12439: out = 14'h1513;
            14'd12440: out = 14'h1513;
            14'd12441: out = 14'h1512;
            14'd12442: out = 14'h1512;
            14'd12443: out = 14'h1511;
            14'd12444: out = 14'h1511;
            14'd12445: out = 14'h1510;
            14'd12446: out = 14'h1510;
            14'd12447: out = 14'h1510;
            14'd12448: out = 14'h150F;
            14'd12449: out = 14'h150F;
            14'd12450: out = 14'h150E;
            14'd12451: out = 14'h150E;
            14'd12452: out = 14'h150D;
            14'd12453: out = 14'h150D;
            14'd12454: out = 14'h150D;
            14'd12455: out = 14'h150C;
            14'd12456: out = 14'h150C;
            14'd12457: out = 14'h150B;
            14'd12458: out = 14'h150B;
            14'd12459: out = 14'h150A;
            14'd12460: out = 14'h150A;
            14'd12461: out = 14'h150A;
            14'd12462: out = 14'h1509;
            14'd12463: out = 14'h1509;
            14'd12464: out = 14'h1508;
            14'd12465: out = 14'h1508;
            14'd12466: out = 14'h1507;
            14'd12467: out = 14'h1507;
            14'd12468: out = 14'h1506;
            14'd12469: out = 14'h1506;
            14'd12470: out = 14'h1506;
            14'd12471: out = 14'h1505;
            14'd12472: out = 14'h1505;
            14'd12473: out = 14'h1504;
            14'd12474: out = 14'h1504;
            14'd12475: out = 14'h1503;
            14'd12476: out = 14'h1503;
            14'd12477: out = 14'h1503;
            14'd12478: out = 14'h1502;
            14'd12479: out = 14'h1502;
            14'd12480: out = 14'h1501;
            14'd12481: out = 14'h1501;
            14'd12482: out = 14'h1500;
            14'd12483: out = 14'h1500;
            14'd12484: out = 14'h1500;
            14'd12485: out = 14'h14FF;
            14'd12486: out = 14'h14FF;
            14'd12487: out = 14'h14FE;
            14'd12488: out = 14'h14FE;
            14'd12489: out = 14'h14FD;
            14'd12490: out = 14'h14FD;
            14'd12491: out = 14'h14FD;
            14'd12492: out = 14'h14FC;
            14'd12493: out = 14'h14FC;
            14'd12494: out = 14'h14FB;
            14'd12495: out = 14'h14FB;
            14'd12496: out = 14'h14FA;
            14'd12497: out = 14'h14FA;
            14'd12498: out = 14'h14FA;
            14'd12499: out = 14'h14F9;
            14'd12500: out = 14'h14F9;
            14'd12501: out = 14'h14F8;
            14'd12502: out = 14'h14F8;
            14'd12503: out = 14'h14F7;
            14'd12504: out = 14'h14F7;
            14'd12505: out = 14'h14F7;
            14'd12506: out = 14'h14F6;
            14'd12507: out = 14'h14F6;
            14'd12508: out = 14'h14F5;
            14'd12509: out = 14'h14F5;
            14'd12510: out = 14'h14F4;
            14'd12511: out = 14'h14F4;
            14'd12512: out = 14'h14F4;
            14'd12513: out = 14'h14F3;
            14'd12514: out = 14'h14F3;
            14'd12515: out = 14'h14F2;
            14'd12516: out = 14'h14F2;
            14'd12517: out = 14'h14F1;
            14'd12518: out = 14'h14F1;
            14'd12519: out = 14'h14F1;
            14'd12520: out = 14'h14F0;
            14'd12521: out = 14'h14F0;
            14'd12522: out = 14'h14EF;
            14'd12523: out = 14'h14EF;
            14'd12524: out = 14'h14EE;
            14'd12525: out = 14'h14EE;
            14'd12526: out = 14'h14EE;
            14'd12527: out = 14'h14ED;
            14'd12528: out = 14'h14ED;
            14'd12529: out = 14'h14EC;
            14'd12530: out = 14'h14EC;
            14'd12531: out = 14'h14EB;
            14'd12532: out = 14'h14EB;
            14'd12533: out = 14'h14EB;
            14'd12534: out = 14'h14EA;
            14'd12535: out = 14'h14EA;
            14'd12536: out = 14'h14E9;
            14'd12537: out = 14'h14E9;
            14'd12538: out = 14'h14E8;
            14'd12539: out = 14'h14E8;
            14'd12540: out = 14'h14E8;
            14'd12541: out = 14'h14E7;
            14'd12542: out = 14'h14E7;
            14'd12543: out = 14'h14E6;
            14'd12544: out = 14'h14E6;
            14'd12545: out = 14'h14E5;
            14'd12546: out = 14'h14E5;
            14'd12547: out = 14'h14E5;
            14'd12548: out = 14'h14E4;
            14'd12549: out = 14'h14E4;
            14'd12550: out = 14'h14E3;
            14'd12551: out = 14'h14E3;
            14'd12552: out = 14'h14E2;
            14'd12553: out = 14'h14E2;
            14'd12554: out = 14'h14E2;
            14'd12555: out = 14'h14E1;
            14'd12556: out = 14'h14E1;
            14'd12557: out = 14'h14E0;
            14'd12558: out = 14'h14E0;
            14'd12559: out = 14'h14DF;
            14'd12560: out = 14'h14DF;
            14'd12561: out = 14'h14DF;
            14'd12562: out = 14'h14DE;
            14'd12563: out = 14'h14DE;
            14'd12564: out = 14'h14DD;
            14'd12565: out = 14'h14DD;
            14'd12566: out = 14'h14DD;
            14'd12567: out = 14'h14DC;
            14'd12568: out = 14'h14DC;
            14'd12569: out = 14'h14DB;
            14'd12570: out = 14'h14DB;
            14'd12571: out = 14'h14DA;
            14'd12572: out = 14'h14DA;
            14'd12573: out = 14'h14DA;
            14'd12574: out = 14'h14D9;
            14'd12575: out = 14'h14D9;
            14'd12576: out = 14'h14D8;
            14'd12577: out = 14'h14D8;
            14'd12578: out = 14'h14D7;
            14'd12579: out = 14'h14D7;
            14'd12580: out = 14'h14D7;
            14'd12581: out = 14'h14D6;
            14'd12582: out = 14'h14D6;
            14'd12583: out = 14'h14D5;
            14'd12584: out = 14'h14D5;
            14'd12585: out = 14'h14D4;
            14'd12586: out = 14'h14D4;
            14'd12587: out = 14'h14D4;
            14'd12588: out = 14'h14D3;
            14'd12589: out = 14'h14D3;
            14'd12590: out = 14'h14D2;
            14'd12591: out = 14'h14D2;
            14'd12592: out = 14'h14D1;
            14'd12593: out = 14'h14D1;
            14'd12594: out = 14'h14D1;
            14'd12595: out = 14'h14D0;
            14'd12596: out = 14'h14D0;
            14'd12597: out = 14'h14CF;
            14'd12598: out = 14'h14CF;
            14'd12599: out = 14'h14CF;
            14'd12600: out = 14'h14CE;
            14'd12601: out = 14'h14CE;
            14'd12602: out = 14'h14CD;
            14'd12603: out = 14'h14CD;
            14'd12604: out = 14'h14CC;
            14'd12605: out = 14'h14CC;
            14'd12606: out = 14'h14CC;
            14'd12607: out = 14'h14CB;
            14'd12608: out = 14'h14CB;
            14'd12609: out = 14'h14CA;
            14'd12610: out = 14'h14CA;
            14'd12611: out = 14'h14C9;
            14'd12612: out = 14'h14C9;
            14'd12613: out = 14'h14C9;
            14'd12614: out = 14'h14C8;
            14'd12615: out = 14'h14C8;
            14'd12616: out = 14'h14C7;
            14'd12617: out = 14'h14C7;
            14'd12618: out = 14'h14C7;
            14'd12619: out = 14'h14C6;
            14'd12620: out = 14'h14C6;
            14'd12621: out = 14'h14C5;
            14'd12622: out = 14'h14C5;
            14'd12623: out = 14'h14C4;
            14'd12624: out = 14'h14C4;
            14'd12625: out = 14'h14C4;
            14'd12626: out = 14'h14C3;
            14'd12627: out = 14'h14C3;
            14'd12628: out = 14'h14C2;
            14'd12629: out = 14'h14C2;
            14'd12630: out = 14'h14C1;
            14'd12631: out = 14'h14C1;
            14'd12632: out = 14'h14C1;
            14'd12633: out = 14'h14C0;
            14'd12634: out = 14'h14C0;
            14'd12635: out = 14'h14BF;
            14'd12636: out = 14'h14BF;
            14'd12637: out = 14'h14BF;
            14'd12638: out = 14'h14BE;
            14'd12639: out = 14'h14BE;
            14'd12640: out = 14'h14BD;
            14'd12641: out = 14'h14BD;
            14'd12642: out = 14'h14BC;
            14'd12643: out = 14'h14BC;
            14'd12644: out = 14'h14BC;
            14'd12645: out = 14'h14BB;
            14'd12646: out = 14'h14BB;
            14'd12647: out = 14'h14BA;
            14'd12648: out = 14'h14BA;
            14'd12649: out = 14'h14B9;
            14'd12650: out = 14'h14B9;
            14'd12651: out = 14'h14B9;
            14'd12652: out = 14'h14B8;
            14'd12653: out = 14'h14B8;
            14'd12654: out = 14'h14B7;
            14'd12655: out = 14'h14B7;
            14'd12656: out = 14'h14B7;
            14'd12657: out = 14'h14B6;
            14'd12658: out = 14'h14B6;
            14'd12659: out = 14'h14B5;
            14'd12660: out = 14'h14B5;
            14'd12661: out = 14'h14B4;
            14'd12662: out = 14'h14B4;
            14'd12663: out = 14'h14B4;
            14'd12664: out = 14'h14B3;
            14'd12665: out = 14'h14B3;
            14'd12666: out = 14'h14B2;
            14'd12667: out = 14'h14B2;
            14'd12668: out = 14'h14B2;
            14'd12669: out = 14'h14B1;
            14'd12670: out = 14'h14B1;
            14'd12671: out = 14'h14B0;
            14'd12672: out = 14'h14B0;
            14'd12673: out = 14'h14AF;
            14'd12674: out = 14'h14AF;
            14'd12675: out = 14'h14AF;
            14'd12676: out = 14'h14AE;
            14'd12677: out = 14'h14AE;
            14'd12678: out = 14'h14AD;
            14'd12679: out = 14'h14AD;
            14'd12680: out = 14'h14AC;
            14'd12681: out = 14'h14AC;
            14'd12682: out = 14'h14AC;
            14'd12683: out = 14'h14AB;
            14'd12684: out = 14'h14AB;
            14'd12685: out = 14'h14AA;
            14'd12686: out = 14'h14AA;
            14'd12687: out = 14'h14AA;
            14'd12688: out = 14'h14A9;
            14'd12689: out = 14'h14A9;
            14'd12690: out = 14'h14A8;
            14'd12691: out = 14'h14A8;
            14'd12692: out = 14'h14A7;
            14'd12693: out = 14'h14A7;
            14'd12694: out = 14'h14A7;
            14'd12695: out = 14'h14A6;
            14'd12696: out = 14'h14A6;
            14'd12697: out = 14'h14A5;
            14'd12698: out = 14'h14A5;
            14'd12699: out = 14'h14A5;
            14'd12700: out = 14'h14A4;
            14'd12701: out = 14'h14A4;
            14'd12702: out = 14'h14A3;
            14'd12703: out = 14'h14A3;
            14'd12704: out = 14'h14A2;
            14'd12705: out = 14'h14A2;
            14'd12706: out = 14'h14A2;
            14'd12707: out = 14'h14A1;
            14'd12708: out = 14'h14A1;
            14'd12709: out = 14'h14A0;
            14'd12710: out = 14'h14A0;
            14'd12711: out = 14'h14A0;
            14'd12712: out = 14'h149F;
            14'd12713: out = 14'h149F;
            14'd12714: out = 14'h149E;
            14'd12715: out = 14'h149E;
            14'd12716: out = 14'h149E;
            14'd12717: out = 14'h149D;
            14'd12718: out = 14'h149D;
            14'd12719: out = 14'h149C;
            14'd12720: out = 14'h149C;
            14'd12721: out = 14'h149B;
            14'd12722: out = 14'h149B;
            14'd12723: out = 14'h149B;
            14'd12724: out = 14'h149A;
            14'd12725: out = 14'h149A;
            14'd12726: out = 14'h1499;
            14'd12727: out = 14'h1499;
            14'd12728: out = 14'h1499;
            14'd12729: out = 14'h1498;
            14'd12730: out = 14'h1498;
            14'd12731: out = 14'h1497;
            14'd12732: out = 14'h1497;
            14'd12733: out = 14'h1496;
            14'd12734: out = 14'h1496;
            14'd12735: out = 14'h1496;
            14'd12736: out = 14'h1495;
            14'd12737: out = 14'h1495;
            14'd12738: out = 14'h1494;
            14'd12739: out = 14'h1494;
            14'd12740: out = 14'h1494;
            14'd12741: out = 14'h1493;
            14'd12742: out = 14'h1493;
            14'd12743: out = 14'h1492;
            14'd12744: out = 14'h1492;
            14'd12745: out = 14'h1492;
            14'd12746: out = 14'h1491;
            14'd12747: out = 14'h1491;
            14'd12748: out = 14'h1490;
            14'd12749: out = 14'h1490;
            14'd12750: out = 14'h148F;
            14'd12751: out = 14'h148F;
            14'd12752: out = 14'h148F;
            14'd12753: out = 14'h148E;
            14'd12754: out = 14'h148E;
            14'd12755: out = 14'h148D;
            14'd12756: out = 14'h148D;
            14'd12757: out = 14'h148D;
            14'd12758: out = 14'h148C;
            14'd12759: out = 14'h148C;
            14'd12760: out = 14'h148B;
            14'd12761: out = 14'h148B;
            14'd12762: out = 14'h148A;
            14'd12763: out = 14'h148A;
            14'd12764: out = 14'h148A;
            14'd12765: out = 14'h1489;
            14'd12766: out = 14'h1489;
            14'd12767: out = 14'h1488;
            14'd12768: out = 14'h1488;
            14'd12769: out = 14'h1488;
            14'd12770: out = 14'h1487;
            14'd12771: out = 14'h1487;
            14'd12772: out = 14'h1486;
            14'd12773: out = 14'h1486;
            14'd12774: out = 14'h1486;
            14'd12775: out = 14'h1485;
            14'd12776: out = 14'h1485;
            14'd12777: out = 14'h1484;
            14'd12778: out = 14'h1484;
            14'd12779: out = 14'h1483;
            14'd12780: out = 14'h1483;
            14'd12781: out = 14'h1483;
            14'd12782: out = 14'h1482;
            14'd12783: out = 14'h1482;
            14'd12784: out = 14'h1481;
            14'd12785: out = 14'h1481;
            14'd12786: out = 14'h1481;
            14'd12787: out = 14'h1480;
            14'd12788: out = 14'h1480;
            14'd12789: out = 14'h147F;
            14'd12790: out = 14'h147F;
            14'd12791: out = 14'h147F;
            14'd12792: out = 14'h147E;
            14'd12793: out = 14'h147E;
            14'd12794: out = 14'h147D;
            14'd12795: out = 14'h147D;
            14'd12796: out = 14'h147D;
            14'd12797: out = 14'h147C;
            14'd12798: out = 14'h147C;
            14'd12799: out = 14'h147B;
            14'd12800: out = 14'h147B;
            14'd12801: out = 14'h147A;
            14'd12802: out = 14'h147A;
            14'd12803: out = 14'h147A;
            14'd12804: out = 14'h1479;
            14'd12805: out = 14'h1479;
            14'd12806: out = 14'h1478;
            14'd12807: out = 14'h1478;
            14'd12808: out = 14'h1478;
            14'd12809: out = 14'h1477;
            14'd12810: out = 14'h1477;
            14'd12811: out = 14'h1476;
            14'd12812: out = 14'h1476;
            14'd12813: out = 14'h1476;
            14'd12814: out = 14'h1475;
            14'd12815: out = 14'h1475;
            14'd12816: out = 14'h1474;
            14'd12817: out = 14'h1474;
            14'd12818: out = 14'h1474;
            14'd12819: out = 14'h1473;
            14'd12820: out = 14'h1473;
            14'd12821: out = 14'h1472;
            14'd12822: out = 14'h1472;
            14'd12823: out = 14'h1471;
            14'd12824: out = 14'h1471;
            14'd12825: out = 14'h1471;
            14'd12826: out = 14'h1470;
            14'd12827: out = 14'h1470;
            14'd12828: out = 14'h146F;
            14'd12829: out = 14'h146F;
            14'd12830: out = 14'h146F;
            14'd12831: out = 14'h146E;
            14'd12832: out = 14'h146E;
            14'd12833: out = 14'h146D;
            14'd12834: out = 14'h146D;
            14'd12835: out = 14'h146D;
            14'd12836: out = 14'h146C;
            14'd12837: out = 14'h146C;
            14'd12838: out = 14'h146B;
            14'd12839: out = 14'h146B;
            14'd12840: out = 14'h146B;
            14'd12841: out = 14'h146A;
            14'd12842: out = 14'h146A;
            14'd12843: out = 14'h1469;
            14'd12844: out = 14'h1469;
            14'd12845: out = 14'h1469;
            14'd12846: out = 14'h1468;
            14'd12847: out = 14'h1468;
            14'd12848: out = 14'h1467;
            14'd12849: out = 14'h1467;
            14'd12850: out = 14'h1466;
            14'd12851: out = 14'h1466;
            14'd12852: out = 14'h1466;
            14'd12853: out = 14'h1465;
            14'd12854: out = 14'h1465;
            14'd12855: out = 14'h1464;
            14'd12856: out = 14'h1464;
            14'd12857: out = 14'h1464;
            14'd12858: out = 14'h1463;
            14'd12859: out = 14'h1463;
            14'd12860: out = 14'h1462;
            14'd12861: out = 14'h1462;
            14'd12862: out = 14'h1462;
            14'd12863: out = 14'h1461;
            14'd12864: out = 14'h1461;
            14'd12865: out = 14'h1460;
            14'd12866: out = 14'h1460;
            14'd12867: out = 14'h1460;
            14'd12868: out = 14'h145F;
            14'd12869: out = 14'h145F;
            14'd12870: out = 14'h145E;
            14'd12871: out = 14'h145E;
            14'd12872: out = 14'h145E;
            14'd12873: out = 14'h145D;
            14'd12874: out = 14'h145D;
            14'd12875: out = 14'h145C;
            14'd12876: out = 14'h145C;
            14'd12877: out = 14'h145C;
            14'd12878: out = 14'h145B;
            14'd12879: out = 14'h145B;
            14'd12880: out = 14'h145A;
            14'd12881: out = 14'h145A;
            14'd12882: out = 14'h145A;
            14'd12883: out = 14'h1459;
            14'd12884: out = 14'h1459;
            14'd12885: out = 14'h1458;
            14'd12886: out = 14'h1458;
            14'd12887: out = 14'h1457;
            14'd12888: out = 14'h1457;
            14'd12889: out = 14'h1457;
            14'd12890: out = 14'h1456;
            14'd12891: out = 14'h1456;
            14'd12892: out = 14'h1455;
            14'd12893: out = 14'h1455;
            14'd12894: out = 14'h1455;
            14'd12895: out = 14'h1454;
            14'd12896: out = 14'h1454;
            14'd12897: out = 14'h1453;
            14'd12898: out = 14'h1453;
            14'd12899: out = 14'h1453;
            14'd12900: out = 14'h1452;
            14'd12901: out = 14'h1452;
            14'd12902: out = 14'h1451;
            14'd12903: out = 14'h1451;
            14'd12904: out = 14'h1451;
            14'd12905: out = 14'h1450;
            14'd12906: out = 14'h1450;
            14'd12907: out = 14'h144F;
            14'd12908: out = 14'h144F;
            14'd12909: out = 14'h144F;
            14'd12910: out = 14'h144E;
            14'd12911: out = 14'h144E;
            14'd12912: out = 14'h144D;
            14'd12913: out = 14'h144D;
            14'd12914: out = 14'h144D;
            14'd12915: out = 14'h144C;
            14'd12916: out = 14'h144C;
            14'd12917: out = 14'h144B;
            14'd12918: out = 14'h144B;
            14'd12919: out = 14'h144B;
            14'd12920: out = 14'h144A;
            14'd12921: out = 14'h144A;
            14'd12922: out = 14'h1449;
            14'd12923: out = 14'h1449;
            14'd12924: out = 14'h1449;
            14'd12925: out = 14'h1448;
            14'd12926: out = 14'h1448;
            14'd12927: out = 14'h1447;
            14'd12928: out = 14'h1447;
            14'd12929: out = 14'h1447;
            14'd12930: out = 14'h1446;
            14'd12931: out = 14'h1446;
            14'd12932: out = 14'h1445;
            14'd12933: out = 14'h1445;
            14'd12934: out = 14'h1445;
            14'd12935: out = 14'h1444;
            14'd12936: out = 14'h1444;
            14'd12937: out = 14'h1443;
            14'd12938: out = 14'h1443;
            14'd12939: out = 14'h1443;
            14'd12940: out = 14'h1442;
            14'd12941: out = 14'h1442;
            14'd12942: out = 14'h1441;
            14'd12943: out = 14'h1441;
            14'd12944: out = 14'h1441;
            14'd12945: out = 14'h1440;
            14'd12946: out = 14'h1440;
            14'd12947: out = 14'h143F;
            14'd12948: out = 14'h143F;
            14'd12949: out = 14'h143F;
            14'd12950: out = 14'h143E;
            14'd12951: out = 14'h143E;
            14'd12952: out = 14'h143D;
            14'd12953: out = 14'h143D;
            14'd12954: out = 14'h143D;
            14'd12955: out = 14'h143C;
            14'd12956: out = 14'h143C;
            14'd12957: out = 14'h143B;
            14'd12958: out = 14'h143B;
            14'd12959: out = 14'h143B;
            14'd12960: out = 14'h143A;
            14'd12961: out = 14'h143A;
            14'd12962: out = 14'h1439;
            14'd12963: out = 14'h1439;
            14'd12964: out = 14'h1439;
            14'd12965: out = 14'h1438;
            14'd12966: out = 14'h1438;
            14'd12967: out = 14'h1437;
            14'd12968: out = 14'h1437;
            14'd12969: out = 14'h1437;
            14'd12970: out = 14'h1436;
            14'd12971: out = 14'h1436;
            14'd12972: out = 14'h1435;
            14'd12973: out = 14'h1435;
            14'd12974: out = 14'h1435;
            14'd12975: out = 14'h1434;
            14'd12976: out = 14'h1434;
            14'd12977: out = 14'h1433;
            14'd12978: out = 14'h1433;
            14'd12979: out = 14'h1433;
            14'd12980: out = 14'h1432;
            14'd12981: out = 14'h1432;
            14'd12982: out = 14'h1431;
            14'd12983: out = 14'h1431;
            14'd12984: out = 14'h1431;
            14'd12985: out = 14'h1430;
            14'd12986: out = 14'h1430;
            14'd12987: out = 14'h142F;
            14'd12988: out = 14'h142F;
            14'd12989: out = 14'h142F;
            14'd12990: out = 14'h142E;
            14'd12991: out = 14'h142E;
            14'd12992: out = 14'h142D;
            14'd12993: out = 14'h142D;
            14'd12994: out = 14'h142D;
            14'd12995: out = 14'h142C;
            14'd12996: out = 14'h142C;
            14'd12997: out = 14'h142B;
            14'd12998: out = 14'h142B;
            14'd12999: out = 14'h142B;
            14'd13000: out = 14'h142A;
            14'd13001: out = 14'h142A;
            14'd13002: out = 14'h1429;
            14'd13003: out = 14'h1429;
            14'd13004: out = 14'h1429;
            14'd13005: out = 14'h1428;
            14'd13006: out = 14'h1428;
            14'd13007: out = 14'h1427;
            14'd13008: out = 14'h1427;
            14'd13009: out = 14'h1427;
            14'd13010: out = 14'h1426;
            14'd13011: out = 14'h1426;
            14'd13012: out = 14'h1425;
            14'd13013: out = 14'h1425;
            14'd13014: out = 14'h1425;
            14'd13015: out = 14'h1424;
            14'd13016: out = 14'h1424;
            14'd13017: out = 14'h1423;
            14'd13018: out = 14'h1423;
            14'd13019: out = 14'h1423;
            14'd13020: out = 14'h1422;
            14'd13021: out = 14'h1422;
            14'd13022: out = 14'h1421;
            14'd13023: out = 14'h1421;
            14'd13024: out = 14'h1421;
            14'd13025: out = 14'h1420;
            14'd13026: out = 14'h1420;
            14'd13027: out = 14'h1420;
            14'd13028: out = 14'h141F;
            14'd13029: out = 14'h141F;
            14'd13030: out = 14'h141E;
            14'd13031: out = 14'h141E;
            14'd13032: out = 14'h141E;
            14'd13033: out = 14'h141D;
            14'd13034: out = 14'h141D;
            14'd13035: out = 14'h141C;
            14'd13036: out = 14'h141C;
            14'd13037: out = 14'h141C;
            14'd13038: out = 14'h141B;
            14'd13039: out = 14'h141B;
            14'd13040: out = 14'h141A;
            14'd13041: out = 14'h141A;
            14'd13042: out = 14'h141A;
            14'd13043: out = 14'h1419;
            14'd13044: out = 14'h1419;
            14'd13045: out = 14'h1418;
            14'd13046: out = 14'h1418;
            14'd13047: out = 14'h1418;
            14'd13048: out = 14'h1417;
            14'd13049: out = 14'h1417;
            14'd13050: out = 14'h1416;
            14'd13051: out = 14'h1416;
            14'd13052: out = 14'h1416;
            14'd13053: out = 14'h1415;
            14'd13054: out = 14'h1415;
            14'd13055: out = 14'h1414;
            14'd13056: out = 14'h1414;
            14'd13057: out = 14'h1414;
            14'd13058: out = 14'h1413;
            14'd13059: out = 14'h1413;
            14'd13060: out = 14'h1413;
            14'd13061: out = 14'h1412;
            14'd13062: out = 14'h1412;
            14'd13063: out = 14'h1411;
            14'd13064: out = 14'h1411;
            14'd13065: out = 14'h1411;
            14'd13066: out = 14'h1410;
            14'd13067: out = 14'h1410;
            14'd13068: out = 14'h140F;
            14'd13069: out = 14'h140F;
            14'd13070: out = 14'h140F;
            14'd13071: out = 14'h140E;
            14'd13072: out = 14'h140E;
            14'd13073: out = 14'h140D;
            14'd13074: out = 14'h140D;
            14'd13075: out = 14'h140D;
            14'd13076: out = 14'h140C;
            14'd13077: out = 14'h140C;
            14'd13078: out = 14'h140B;
            14'd13079: out = 14'h140B;
            14'd13080: out = 14'h140B;
            14'd13081: out = 14'h140A;
            14'd13082: out = 14'h140A;
            14'd13083: out = 14'h1409;
            14'd13084: out = 14'h1409;
            14'd13085: out = 14'h1409;
            14'd13086: out = 14'h1408;
            14'd13087: out = 14'h1408;
            14'd13088: out = 14'h1408;
            14'd13089: out = 14'h1407;
            14'd13090: out = 14'h1407;
            14'd13091: out = 14'h1406;
            14'd13092: out = 14'h1406;
            14'd13093: out = 14'h1406;
            14'd13094: out = 14'h1405;
            14'd13095: out = 14'h1405;
            14'd13096: out = 14'h1404;
            14'd13097: out = 14'h1404;
            14'd13098: out = 14'h1404;
            14'd13099: out = 14'h1403;
            14'd13100: out = 14'h1403;
            14'd13101: out = 14'h1402;
            14'd13102: out = 14'h1402;
            14'd13103: out = 14'h1402;
            14'd13104: out = 14'h1401;
            14'd13105: out = 14'h1401;
            14'd13106: out = 14'h1400;
            14'd13107: out = 14'h1400;
            14'd13108: out = 14'h1400;
            14'd13109: out = 14'h13FF;
            14'd13110: out = 14'h13FF;
            14'd13111: out = 14'h13FF;
            14'd13112: out = 14'h13FE;
            14'd13113: out = 14'h13FE;
            14'd13114: out = 14'h13FD;
            14'd13115: out = 14'h13FD;
            14'd13116: out = 14'h13FD;
            14'd13117: out = 14'h13FC;
            14'd13118: out = 14'h13FC;
            14'd13119: out = 14'h13FB;
            14'd13120: out = 14'h13FB;
            14'd13121: out = 14'h13FB;
            14'd13122: out = 14'h13FA;
            14'd13123: out = 14'h13FA;
            14'd13124: out = 14'h13F9;
            14'd13125: out = 14'h13F9;
            14'd13126: out = 14'h13F9;
            14'd13127: out = 14'h13F8;
            14'd13128: out = 14'h13F8;
            14'd13129: out = 14'h13F7;
            14'd13130: out = 14'h13F7;
            14'd13131: out = 14'h13F7;
            14'd13132: out = 14'h13F6;
            14'd13133: out = 14'h13F6;
            14'd13134: out = 14'h13F6;
            14'd13135: out = 14'h13F5;
            14'd13136: out = 14'h13F5;
            14'd13137: out = 14'h13F4;
            14'd13138: out = 14'h13F4;
            14'd13139: out = 14'h13F4;
            14'd13140: out = 14'h13F3;
            14'd13141: out = 14'h13F3;
            14'd13142: out = 14'h13F2;
            14'd13143: out = 14'h13F2;
            14'd13144: out = 14'h13F2;
            14'd13145: out = 14'h13F1;
            14'd13146: out = 14'h13F1;
            14'd13147: out = 14'h13F1;
            14'd13148: out = 14'h13F0;
            14'd13149: out = 14'h13F0;
            14'd13150: out = 14'h13EF;
            14'd13151: out = 14'h13EF;
            14'd13152: out = 14'h13EF;
            14'd13153: out = 14'h13EE;
            14'd13154: out = 14'h13EE;
            14'd13155: out = 14'h13ED;
            14'd13156: out = 14'h13ED;
            14'd13157: out = 14'h13ED;
            14'd13158: out = 14'h13EC;
            14'd13159: out = 14'h13EC;
            14'd13160: out = 14'h13EB;
            14'd13161: out = 14'h13EB;
            14'd13162: out = 14'h13EB;
            14'd13163: out = 14'h13EA;
            14'd13164: out = 14'h13EA;
            14'd13165: out = 14'h13EA;
            14'd13166: out = 14'h13E9;
            14'd13167: out = 14'h13E9;
            14'd13168: out = 14'h13E8;
            14'd13169: out = 14'h13E8;
            14'd13170: out = 14'h13E8;
            14'd13171: out = 14'h13E7;
            14'd13172: out = 14'h13E7;
            14'd13173: out = 14'h13E6;
            14'd13174: out = 14'h13E6;
            14'd13175: out = 14'h13E6;
            14'd13176: out = 14'h13E5;
            14'd13177: out = 14'h13E5;
            14'd13178: out = 14'h13E4;
            14'd13179: out = 14'h13E4;
            14'd13180: out = 14'h13E4;
            14'd13181: out = 14'h13E3;
            14'd13182: out = 14'h13E3;
            14'd13183: out = 14'h13E3;
            14'd13184: out = 14'h13E2;
            14'd13185: out = 14'h13E2;
            14'd13186: out = 14'h13E1;
            14'd13187: out = 14'h13E1;
            14'd13188: out = 14'h13E1;
            14'd13189: out = 14'h13E0;
            14'd13190: out = 14'h13E0;
            14'd13191: out = 14'h13DF;
            14'd13192: out = 14'h13DF;
            14'd13193: out = 14'h13DF;
            14'd13194: out = 14'h13DE;
            14'd13195: out = 14'h13DE;
            14'd13196: out = 14'h13DE;
            14'd13197: out = 14'h13DD;
            14'd13198: out = 14'h13DD;
            14'd13199: out = 14'h13DC;
            14'd13200: out = 14'h13DC;
            14'd13201: out = 14'h13DC;
            14'd13202: out = 14'h13DB;
            14'd13203: out = 14'h13DB;
            14'd13204: out = 14'h13DA;
            14'd13205: out = 14'h13DA;
            14'd13206: out = 14'h13DA;
            14'd13207: out = 14'h13D9;
            14'd13208: out = 14'h13D9;
            14'd13209: out = 14'h13D9;
            14'd13210: out = 14'h13D8;
            14'd13211: out = 14'h13D8;
            14'd13212: out = 14'h13D7;
            14'd13213: out = 14'h13D7;
            14'd13214: out = 14'h13D7;
            14'd13215: out = 14'h13D6;
            14'd13216: out = 14'h13D6;
            14'd13217: out = 14'h13D5;
            14'd13218: out = 14'h13D5;
            14'd13219: out = 14'h13D5;
            14'd13220: out = 14'h13D4;
            14'd13221: out = 14'h13D4;
            14'd13222: out = 14'h13D4;
            14'd13223: out = 14'h13D3;
            14'd13224: out = 14'h13D3;
            14'd13225: out = 14'h13D2;
            14'd13226: out = 14'h13D2;
            14'd13227: out = 14'h13D2;
            14'd13228: out = 14'h13D1;
            14'd13229: out = 14'h13D1;
            14'd13230: out = 14'h13D0;
            14'd13231: out = 14'h13D0;
            14'd13232: out = 14'h13D0;
            14'd13233: out = 14'h13CF;
            14'd13234: out = 14'h13CF;
            14'd13235: out = 14'h13CF;
            14'd13236: out = 14'h13CE;
            14'd13237: out = 14'h13CE;
            14'd13238: out = 14'h13CD;
            14'd13239: out = 14'h13CD;
            14'd13240: out = 14'h13CD;
            14'd13241: out = 14'h13CC;
            14'd13242: out = 14'h13CC;
            14'd13243: out = 14'h13CB;
            14'd13244: out = 14'h13CB;
            14'd13245: out = 14'h13CB;
            14'd13246: out = 14'h13CA;
            14'd13247: out = 14'h13CA;
            14'd13248: out = 14'h13CA;
            14'd13249: out = 14'h13C9;
            14'd13250: out = 14'h13C9;
            14'd13251: out = 14'h13C8;
            14'd13252: out = 14'h13C8;
            14'd13253: out = 14'h13C8;
            14'd13254: out = 14'h13C7;
            14'd13255: out = 14'h13C7;
            14'd13256: out = 14'h13C7;
            14'd13257: out = 14'h13C6;
            14'd13258: out = 14'h13C6;
            14'd13259: out = 14'h13C5;
            14'd13260: out = 14'h13C5;
            14'd13261: out = 14'h13C5;
            14'd13262: out = 14'h13C4;
            14'd13263: out = 14'h13C4;
            14'd13264: out = 14'h13C3;
            14'd13265: out = 14'h13C3;
            14'd13266: out = 14'h13C3;
            14'd13267: out = 14'h13C2;
            14'd13268: out = 14'h13C2;
            14'd13269: out = 14'h13C2;
            14'd13270: out = 14'h13C1;
            14'd13271: out = 14'h13C1;
            14'd13272: out = 14'h13C0;
            14'd13273: out = 14'h13C0;
            14'd13274: out = 14'h13C0;
            14'd13275: out = 14'h13BF;
            14'd13276: out = 14'h13BF;
            14'd13277: out = 14'h13BF;
            14'd13278: out = 14'h13BE;
            14'd13279: out = 14'h13BE;
            14'd13280: out = 14'h13BD;
            14'd13281: out = 14'h13BD;
            14'd13282: out = 14'h13BD;
            14'd13283: out = 14'h13BC;
            14'd13284: out = 14'h13BC;
            14'd13285: out = 14'h13BB;
            14'd13286: out = 14'h13BB;
            14'd13287: out = 14'h13BB;
            14'd13288: out = 14'h13BA;
            14'd13289: out = 14'h13BA;
            14'd13290: out = 14'h13BA;
            14'd13291: out = 14'h13B9;
            14'd13292: out = 14'h13B9;
            14'd13293: out = 14'h13B8;
            14'd13294: out = 14'h13B8;
            14'd13295: out = 14'h13B8;
            14'd13296: out = 14'h13B7;
            14'd13297: out = 14'h13B7;
            14'd13298: out = 14'h13B7;
            14'd13299: out = 14'h13B6;
            14'd13300: out = 14'h13B6;
            14'd13301: out = 14'h13B5;
            14'd13302: out = 14'h13B5;
            14'd13303: out = 14'h13B5;
            14'd13304: out = 14'h13B4;
            14'd13305: out = 14'h13B4;
            14'd13306: out = 14'h13B4;
            14'd13307: out = 14'h13B3;
            14'd13308: out = 14'h13B3;
            14'd13309: out = 14'h13B2;
            14'd13310: out = 14'h13B2;
            14'd13311: out = 14'h13B2;
            14'd13312: out = 14'h13B1;
            14'd13313: out = 14'h13B1;
            14'd13314: out = 14'h13B0;
            14'd13315: out = 14'h13B0;
            14'd13316: out = 14'h13B0;
            14'd13317: out = 14'h13AF;
            14'd13318: out = 14'h13AF;
            14'd13319: out = 14'h13AF;
            14'd13320: out = 14'h13AE;
            14'd13321: out = 14'h13AE;
            14'd13322: out = 14'h13AD;
            14'd13323: out = 14'h13AD;
            14'd13324: out = 14'h13AD;
            14'd13325: out = 14'h13AC;
            14'd13326: out = 14'h13AC;
            14'd13327: out = 14'h13AC;
            14'd13328: out = 14'h13AB;
            14'd13329: out = 14'h13AB;
            14'd13330: out = 14'h13AA;
            14'd13331: out = 14'h13AA;
            14'd13332: out = 14'h13AA;
            14'd13333: out = 14'h13A9;
            14'd13334: out = 14'h13A9;
            14'd13335: out = 14'h13A9;
            14'd13336: out = 14'h13A8;
            14'd13337: out = 14'h13A8;
            14'd13338: out = 14'h13A7;
            14'd13339: out = 14'h13A7;
            14'd13340: out = 14'h13A7;
            14'd13341: out = 14'h13A6;
            14'd13342: out = 14'h13A6;
            14'd13343: out = 14'h13A6;
            14'd13344: out = 14'h13A5;
            14'd13345: out = 14'h13A5;
            14'd13346: out = 14'h13A4;
            14'd13347: out = 14'h13A4;
            14'd13348: out = 14'h13A4;
            14'd13349: out = 14'h13A3;
            14'd13350: out = 14'h13A3;
            14'd13351: out = 14'h13A3;
            14'd13352: out = 14'h13A2;
            14'd13353: out = 14'h13A2;
            14'd13354: out = 14'h13A1;
            14'd13355: out = 14'h13A1;
            14'd13356: out = 14'h13A1;
            14'd13357: out = 14'h13A0;
            14'd13358: out = 14'h13A0;
            14'd13359: out = 14'h139F;
            14'd13360: out = 14'h139F;
            14'd13361: out = 14'h139F;
            14'd13362: out = 14'h139E;
            14'd13363: out = 14'h139E;
            14'd13364: out = 14'h139E;
            14'd13365: out = 14'h139D;
            14'd13366: out = 14'h139D;
            14'd13367: out = 14'h139C;
            14'd13368: out = 14'h139C;
            14'd13369: out = 14'h139C;
            14'd13370: out = 14'h139B;
            14'd13371: out = 14'h139B;
            14'd13372: out = 14'h139B;
            14'd13373: out = 14'h139A;
            14'd13374: out = 14'h139A;
            14'd13375: out = 14'h1399;
            14'd13376: out = 14'h1399;
            14'd13377: out = 14'h1399;
            14'd13378: out = 14'h1398;
            14'd13379: out = 14'h1398;
            14'd13380: out = 14'h1398;
            14'd13381: out = 14'h1397;
            14'd13382: out = 14'h1397;
            14'd13383: out = 14'h1396;
            14'd13384: out = 14'h1396;
            14'd13385: out = 14'h1396;
            14'd13386: out = 14'h1395;
            14'd13387: out = 14'h1395;
            14'd13388: out = 14'h1395;
            14'd13389: out = 14'h1394;
            14'd13390: out = 14'h1394;
            14'd13391: out = 14'h1393;
            14'd13392: out = 14'h1393;
            14'd13393: out = 14'h1393;
            14'd13394: out = 14'h1392;
            14'd13395: out = 14'h1392;
            14'd13396: out = 14'h1392;
            14'd13397: out = 14'h1391;
            14'd13398: out = 14'h1391;
            14'd13399: out = 14'h1390;
            14'd13400: out = 14'h1390;
            14'd13401: out = 14'h1390;
            14'd13402: out = 14'h138F;
            14'd13403: out = 14'h138F;
            14'd13404: out = 14'h138F;
            14'd13405: out = 14'h138E;
            14'd13406: out = 14'h138E;
            14'd13407: out = 14'h138E;
            14'd13408: out = 14'h138D;
            14'd13409: out = 14'h138D;
            14'd13410: out = 14'h138C;
            14'd13411: out = 14'h138C;
            14'd13412: out = 14'h138C;
            14'd13413: out = 14'h138B;
            14'd13414: out = 14'h138B;
            14'd13415: out = 14'h138B;
            14'd13416: out = 14'h138A;
            14'd13417: out = 14'h138A;
            14'd13418: out = 14'h1389;
            14'd13419: out = 14'h1389;
            14'd13420: out = 14'h1389;
            14'd13421: out = 14'h1388;
            14'd13422: out = 14'h1388;
            14'd13423: out = 14'h1388;
            14'd13424: out = 14'h1387;
            14'd13425: out = 14'h1387;
            14'd13426: out = 14'h1386;
            14'd13427: out = 14'h1386;
            14'd13428: out = 14'h1386;
            14'd13429: out = 14'h1385;
            14'd13430: out = 14'h1385;
            14'd13431: out = 14'h1385;
            14'd13432: out = 14'h1384;
            14'd13433: out = 14'h1384;
            14'd13434: out = 14'h1383;
            14'd13435: out = 14'h1383;
            14'd13436: out = 14'h1383;
            14'd13437: out = 14'h1382;
            14'd13438: out = 14'h1382;
            14'd13439: out = 14'h1382;
            14'd13440: out = 14'h1381;
            14'd13441: out = 14'h1381;
            14'd13442: out = 14'h1380;
            14'd13443: out = 14'h1380;
            14'd13444: out = 14'h1380;
            14'd13445: out = 14'h137F;
            14'd13446: out = 14'h137F;
            14'd13447: out = 14'h137F;
            14'd13448: out = 14'h137E;
            14'd13449: out = 14'h137E;
            14'd13450: out = 14'h137E;
            14'd13451: out = 14'h137D;
            14'd13452: out = 14'h137D;
            14'd13453: out = 14'h137C;
            14'd13454: out = 14'h137C;
            14'd13455: out = 14'h137C;
            14'd13456: out = 14'h137B;
            14'd13457: out = 14'h137B;
            14'd13458: out = 14'h137B;
            14'd13459: out = 14'h137A;
            14'd13460: out = 14'h137A;
            14'd13461: out = 14'h1379;
            14'd13462: out = 14'h1379;
            14'd13463: out = 14'h1379;
            14'd13464: out = 14'h1378;
            14'd13465: out = 14'h1378;
            14'd13466: out = 14'h1378;
            14'd13467: out = 14'h1377;
            14'd13468: out = 14'h1377;
            14'd13469: out = 14'h1376;
            14'd13470: out = 14'h1376;
            14'd13471: out = 14'h1376;
            14'd13472: out = 14'h1375;
            14'd13473: out = 14'h1375;
            14'd13474: out = 14'h1375;
            14'd13475: out = 14'h1374;
            14'd13476: out = 14'h1374;
            14'd13477: out = 14'h1374;
            14'd13478: out = 14'h1373;
            14'd13479: out = 14'h1373;
            14'd13480: out = 14'h1372;
            14'd13481: out = 14'h1372;
            14'd13482: out = 14'h1372;
            14'd13483: out = 14'h1371;
            14'd13484: out = 14'h1371;
            14'd13485: out = 14'h1371;
            14'd13486: out = 14'h1370;
            14'd13487: out = 14'h1370;
            14'd13488: out = 14'h136F;
            14'd13489: out = 14'h136F;
            14'd13490: out = 14'h136F;
            14'd13491: out = 14'h136E;
            14'd13492: out = 14'h136E;
            14'd13493: out = 14'h136E;
            14'd13494: out = 14'h136D;
            14'd13495: out = 14'h136D;
            14'd13496: out = 14'h136D;
            14'd13497: out = 14'h136C;
            14'd13498: out = 14'h136C;
            14'd13499: out = 14'h136B;
            14'd13500: out = 14'h136B;
            14'd13501: out = 14'h136B;
            14'd13502: out = 14'h136A;
            14'd13503: out = 14'h136A;
            14'd13504: out = 14'h136A;
            14'd13505: out = 14'h1369;
            14'd13506: out = 14'h1369;
            14'd13507: out = 14'h1368;
            14'd13508: out = 14'h1368;
            14'd13509: out = 14'h1368;
            14'd13510: out = 14'h1367;
            14'd13511: out = 14'h1367;
            14'd13512: out = 14'h1367;
            14'd13513: out = 14'h1366;
            14'd13514: out = 14'h1366;
            14'd13515: out = 14'h1366;
            14'd13516: out = 14'h1365;
            14'd13517: out = 14'h1365;
            14'd13518: out = 14'h1364;
            14'd13519: out = 14'h1364;
            14'd13520: out = 14'h1364;
            14'd13521: out = 14'h1363;
            14'd13522: out = 14'h1363;
            14'd13523: out = 14'h1363;
            14'd13524: out = 14'h1362;
            14'd13525: out = 14'h1362;
            14'd13526: out = 14'h1361;
            14'd13527: out = 14'h1361;
            14'd13528: out = 14'h1361;
            14'd13529: out = 14'h1360;
            14'd13530: out = 14'h1360;
            14'd13531: out = 14'h1360;
            14'd13532: out = 14'h135F;
            14'd13533: out = 14'h135F;
            14'd13534: out = 14'h135F;
            14'd13535: out = 14'h135E;
            14'd13536: out = 14'h135E;
            14'd13537: out = 14'h135D;
            14'd13538: out = 14'h135D;
            14'd13539: out = 14'h135D;
            14'd13540: out = 14'h135C;
            14'd13541: out = 14'h135C;
            14'd13542: out = 14'h135C;
            14'd13543: out = 14'h135B;
            14'd13544: out = 14'h135B;
            14'd13545: out = 14'h135B;
            14'd13546: out = 14'h135A;
            14'd13547: out = 14'h135A;
            14'd13548: out = 14'h1359;
            14'd13549: out = 14'h1359;
            14'd13550: out = 14'h1359;
            14'd13551: out = 14'h1358;
            14'd13552: out = 14'h1358;
            14'd13553: out = 14'h1358;
            14'd13554: out = 14'h1357;
            14'd13555: out = 14'h1357;
            14'd13556: out = 14'h1356;
            14'd13557: out = 14'h1356;
            14'd13558: out = 14'h1356;
            14'd13559: out = 14'h1355;
            14'd13560: out = 14'h1355;
            14'd13561: out = 14'h1355;
            14'd13562: out = 14'h1354;
            14'd13563: out = 14'h1354;
            14'd13564: out = 14'h1354;
            14'd13565: out = 14'h1353;
            14'd13566: out = 14'h1353;
            14'd13567: out = 14'h1352;
            14'd13568: out = 14'h1352;
            14'd13569: out = 14'h1352;
            14'd13570: out = 14'h1351;
            14'd13571: out = 14'h1351;
            14'd13572: out = 14'h1351;
            14'd13573: out = 14'h1350;
            14'd13574: out = 14'h1350;
            14'd13575: out = 14'h1350;
            14'd13576: out = 14'h134F;
            14'd13577: out = 14'h134F;
            14'd13578: out = 14'h134E;
            14'd13579: out = 14'h134E;
            14'd13580: out = 14'h134E;
            14'd13581: out = 14'h134D;
            14'd13582: out = 14'h134D;
            14'd13583: out = 14'h134D;
            14'd13584: out = 14'h134C;
            14'd13585: out = 14'h134C;
            14'd13586: out = 14'h134C;
            14'd13587: out = 14'h134B;
            14'd13588: out = 14'h134B;
            14'd13589: out = 14'h134A;
            14'd13590: out = 14'h134A;
            14'd13591: out = 14'h134A;
            14'd13592: out = 14'h1349;
            14'd13593: out = 14'h1349;
            14'd13594: out = 14'h1349;
            14'd13595: out = 14'h1348;
            14'd13596: out = 14'h1348;
            14'd13597: out = 14'h1348;
            14'd13598: out = 14'h1347;
            14'd13599: out = 14'h1347;
            14'd13600: out = 14'h1346;
            14'd13601: out = 14'h1346;
            14'd13602: out = 14'h1346;
            14'd13603: out = 14'h1345;
            14'd13604: out = 14'h1345;
            14'd13605: out = 14'h1345;
            14'd13606: out = 14'h1344;
            14'd13607: out = 14'h1344;
            14'd13608: out = 14'h1344;
            14'd13609: out = 14'h1343;
            14'd13610: out = 14'h1343;
            14'd13611: out = 14'h1342;
            14'd13612: out = 14'h1342;
            14'd13613: out = 14'h1342;
            14'd13614: out = 14'h1341;
            14'd13615: out = 14'h1341;
            14'd13616: out = 14'h1341;
            14'd13617: out = 14'h1340;
            14'd13618: out = 14'h1340;
            14'd13619: out = 14'h1340;
            14'd13620: out = 14'h133F;
            14'd13621: out = 14'h133F;
            14'd13622: out = 14'h133F;
            14'd13623: out = 14'h133E;
            14'd13624: out = 14'h133E;
            14'd13625: out = 14'h133D;
            14'd13626: out = 14'h133D;
            14'd13627: out = 14'h133D;
            14'd13628: out = 14'h133C;
            14'd13629: out = 14'h133C;
            14'd13630: out = 14'h133C;
            14'd13631: out = 14'h133B;
            14'd13632: out = 14'h133B;
            14'd13633: out = 14'h133B;
            14'd13634: out = 14'h133A;
            14'd13635: out = 14'h133A;
            14'd13636: out = 14'h1339;
            14'd13637: out = 14'h1339;
            14'd13638: out = 14'h1339;
            14'd13639: out = 14'h1338;
            14'd13640: out = 14'h1338;
            14'd13641: out = 14'h1338;
            14'd13642: out = 14'h1337;
            14'd13643: out = 14'h1337;
            14'd13644: out = 14'h1337;
            14'd13645: out = 14'h1336;
            14'd13646: out = 14'h1336;
            14'd13647: out = 14'h1335;
            14'd13648: out = 14'h1335;
            14'd13649: out = 14'h1335;
            14'd13650: out = 14'h1334;
            14'd13651: out = 14'h1334;
            14'd13652: out = 14'h1334;
            14'd13653: out = 14'h1333;
            14'd13654: out = 14'h1333;
            14'd13655: out = 14'h1333;
            14'd13656: out = 14'h1332;
            14'd13657: out = 14'h1332;
            14'd13658: out = 14'h1332;
            14'd13659: out = 14'h1331;
            14'd13660: out = 14'h1331;
            14'd13661: out = 14'h1330;
            14'd13662: out = 14'h1330;
            14'd13663: out = 14'h1330;
            14'd13664: out = 14'h132F;
            14'd13665: out = 14'h132F;
            14'd13666: out = 14'h132F;
            14'd13667: out = 14'h132E;
            14'd13668: out = 14'h132E;
            14'd13669: out = 14'h132E;
            14'd13670: out = 14'h132D;
            14'd13671: out = 14'h132D;
            14'd13672: out = 14'h132C;
            14'd13673: out = 14'h132C;
            14'd13674: out = 14'h132C;
            14'd13675: out = 14'h132B;
            14'd13676: out = 14'h132B;
            14'd13677: out = 14'h132B;
            14'd13678: out = 14'h132A;
            14'd13679: out = 14'h132A;
            14'd13680: out = 14'h132A;
            14'd13681: out = 14'h1329;
            14'd13682: out = 14'h1329;
            14'd13683: out = 14'h1329;
            14'd13684: out = 14'h1328;
            14'd13685: out = 14'h1328;
            14'd13686: out = 14'h1327;
            14'd13687: out = 14'h1327;
            14'd13688: out = 14'h1327;
            14'd13689: out = 14'h1326;
            14'd13690: out = 14'h1326;
            14'd13691: out = 14'h1326;
            14'd13692: out = 14'h1325;
            14'd13693: out = 14'h1325;
            14'd13694: out = 14'h1325;
            14'd13695: out = 14'h1324;
            14'd13696: out = 14'h1324;
            14'd13697: out = 14'h1324;
            14'd13698: out = 14'h1323;
            14'd13699: out = 14'h1323;
            14'd13700: out = 14'h1322;
            14'd13701: out = 14'h1322;
            14'd13702: out = 14'h1322;
            14'd13703: out = 14'h1321;
            14'd13704: out = 14'h1321;
            14'd13705: out = 14'h1321;
            14'd13706: out = 14'h1320;
            14'd13707: out = 14'h1320;
            14'd13708: out = 14'h1320;
            14'd13709: out = 14'h131F;
            14'd13710: out = 14'h131F;
            14'd13711: out = 14'h131F;
            14'd13712: out = 14'h131E;
            14'd13713: out = 14'h131E;
            14'd13714: out = 14'h131D;
            14'd13715: out = 14'h131D;
            14'd13716: out = 14'h131D;
            14'd13717: out = 14'h131C;
            14'd13718: out = 14'h131C;
            14'd13719: out = 14'h131C;
            14'd13720: out = 14'h131B;
            14'd13721: out = 14'h131B;
            14'd13722: out = 14'h131B;
            14'd13723: out = 14'h131A;
            14'd13724: out = 14'h131A;
            14'd13725: out = 14'h131A;
            14'd13726: out = 14'h1319;
            14'd13727: out = 14'h1319;
            14'd13728: out = 14'h1318;
            14'd13729: out = 14'h1318;
            14'd13730: out = 14'h1318;
            14'd13731: out = 14'h1317;
            14'd13732: out = 14'h1317;
            14'd13733: out = 14'h1317;
            14'd13734: out = 14'h1316;
            14'd13735: out = 14'h1316;
            14'd13736: out = 14'h1316;
            14'd13737: out = 14'h1315;
            14'd13738: out = 14'h1315;
            14'd13739: out = 14'h1315;
            14'd13740: out = 14'h1314;
            14'd13741: out = 14'h1314;
            14'd13742: out = 14'h1313;
            14'd13743: out = 14'h1313;
            14'd13744: out = 14'h1313;
            14'd13745: out = 14'h1312;
            14'd13746: out = 14'h1312;
            14'd13747: out = 14'h1312;
            14'd13748: out = 14'h1311;
            14'd13749: out = 14'h1311;
            14'd13750: out = 14'h1311;
            14'd13751: out = 14'h1310;
            14'd13752: out = 14'h1310;
            14'd13753: out = 14'h1310;
            14'd13754: out = 14'h130F;
            14'd13755: out = 14'h130F;
            14'd13756: out = 14'h130F;
            14'd13757: out = 14'h130E;
            14'd13758: out = 14'h130E;
            14'd13759: out = 14'h130D;
            14'd13760: out = 14'h130D;
            14'd13761: out = 14'h130D;
            14'd13762: out = 14'h130C;
            14'd13763: out = 14'h130C;
            14'd13764: out = 14'h130C;
            14'd13765: out = 14'h130B;
            14'd13766: out = 14'h130B;
            14'd13767: out = 14'h130B;
            14'd13768: out = 14'h130A;
            14'd13769: out = 14'h130A;
            14'd13770: out = 14'h130A;
            14'd13771: out = 14'h1309;
            14'd13772: out = 14'h1309;
            14'd13773: out = 14'h1308;
            14'd13774: out = 14'h1308;
            14'd13775: out = 14'h1308;
            14'd13776: out = 14'h1307;
            14'd13777: out = 14'h1307;
            14'd13778: out = 14'h1307;
            14'd13779: out = 14'h1306;
            14'd13780: out = 14'h1306;
            14'd13781: out = 14'h1306;
            14'd13782: out = 14'h1305;
            14'd13783: out = 14'h1305;
            14'd13784: out = 14'h1305;
            14'd13785: out = 14'h1304;
            14'd13786: out = 14'h1304;
            14'd13787: out = 14'h1304;
            14'd13788: out = 14'h1303;
            14'd13789: out = 14'h1303;
            14'd13790: out = 14'h1302;
            14'd13791: out = 14'h1302;
            14'd13792: out = 14'h1302;
            14'd13793: out = 14'h1301;
            14'd13794: out = 14'h1301;
            14'd13795: out = 14'h1301;
            14'd13796: out = 14'h1300;
            14'd13797: out = 14'h1300;
            14'd13798: out = 14'h1300;
            14'd13799: out = 14'h12FF;
            14'd13800: out = 14'h12FF;
            14'd13801: out = 14'h12FF;
            14'd13802: out = 14'h12FE;
            14'd13803: out = 14'h12FE;
            14'd13804: out = 14'h12FE;
            14'd13805: out = 14'h12FD;
            14'd13806: out = 14'h12FD;
            14'd13807: out = 14'h12FC;
            14'd13808: out = 14'h12FC;
            14'd13809: out = 14'h12FC;
            14'd13810: out = 14'h12FB;
            14'd13811: out = 14'h12FB;
            14'd13812: out = 14'h12FB;
            14'd13813: out = 14'h12FA;
            14'd13814: out = 14'h12FA;
            14'd13815: out = 14'h12FA;
            14'd13816: out = 14'h12F9;
            14'd13817: out = 14'h12F9;
            14'd13818: out = 14'h12F9;
            14'd13819: out = 14'h12F8;
            14'd13820: out = 14'h12F8;
            14'd13821: out = 14'h12F8;
            14'd13822: out = 14'h12F7;
            14'd13823: out = 14'h12F7;
            14'd13824: out = 14'h12F7;
            14'd13825: out = 14'h12F6;
            14'd13826: out = 14'h12F6;
            14'd13827: out = 14'h12F5;
            14'd13828: out = 14'h12F5;
            14'd13829: out = 14'h12F5;
            14'd13830: out = 14'h12F4;
            14'd13831: out = 14'h12F4;
            14'd13832: out = 14'h12F4;
            14'd13833: out = 14'h12F3;
            14'd13834: out = 14'h12F3;
            14'd13835: out = 14'h12F3;
            14'd13836: out = 14'h12F2;
            14'd13837: out = 14'h12F2;
            14'd13838: out = 14'h12F2;
            14'd13839: out = 14'h12F1;
            14'd13840: out = 14'h12F1;
            14'd13841: out = 14'h12F1;
            14'd13842: out = 14'h12F0;
            14'd13843: out = 14'h12F0;
            14'd13844: out = 14'h12F0;
            14'd13845: out = 14'h12EF;
            14'd13846: out = 14'h12EF;
            14'd13847: out = 14'h12EE;
            14'd13848: out = 14'h12EE;
            14'd13849: out = 14'h12EE;
            14'd13850: out = 14'h12ED;
            14'd13851: out = 14'h12ED;
            14'd13852: out = 14'h12ED;
            14'd13853: out = 14'h12EC;
            14'd13854: out = 14'h12EC;
            14'd13855: out = 14'h12EC;
            14'd13856: out = 14'h12EB;
            14'd13857: out = 14'h12EB;
            14'd13858: out = 14'h12EB;
            14'd13859: out = 14'h12EA;
            14'd13860: out = 14'h12EA;
            14'd13861: out = 14'h12EA;
            14'd13862: out = 14'h12E9;
            14'd13863: out = 14'h12E9;
            14'd13864: out = 14'h12E9;
            14'd13865: out = 14'h12E8;
            14'd13866: out = 14'h12E8;
            14'd13867: out = 14'h12E7;
            14'd13868: out = 14'h12E7;
            14'd13869: out = 14'h12E7;
            14'd13870: out = 14'h12E6;
            14'd13871: out = 14'h12E6;
            14'd13872: out = 14'h12E6;
            14'd13873: out = 14'h12E5;
            14'd13874: out = 14'h12E5;
            14'd13875: out = 14'h12E5;
            14'd13876: out = 14'h12E4;
            14'd13877: out = 14'h12E4;
            14'd13878: out = 14'h12E4;
            14'd13879: out = 14'h12E3;
            14'd13880: out = 14'h12E3;
            14'd13881: out = 14'h12E3;
            14'd13882: out = 14'h12E2;
            14'd13883: out = 14'h12E2;
            14'd13884: out = 14'h12E2;
            14'd13885: out = 14'h12E1;
            14'd13886: out = 14'h12E1;
            14'd13887: out = 14'h12E0;
            14'd13888: out = 14'h12E0;
            14'd13889: out = 14'h12E0;
            14'd13890: out = 14'h12DF;
            14'd13891: out = 14'h12DF;
            14'd13892: out = 14'h12DF;
            14'd13893: out = 14'h12DE;
            14'd13894: out = 14'h12DE;
            14'd13895: out = 14'h12DE;
            14'd13896: out = 14'h12DD;
            14'd13897: out = 14'h12DD;
            14'd13898: out = 14'h12DD;
            14'd13899: out = 14'h12DC;
            14'd13900: out = 14'h12DC;
            14'd13901: out = 14'h12DC;
            14'd13902: out = 14'h12DB;
            14'd13903: out = 14'h12DB;
            14'd13904: out = 14'h12DB;
            14'd13905: out = 14'h12DA;
            14'd13906: out = 14'h12DA;
            14'd13907: out = 14'h12DA;
            14'd13908: out = 14'h12D9;
            14'd13909: out = 14'h12D9;
            14'd13910: out = 14'h12D9;
            14'd13911: out = 14'h12D8;
            14'd13912: out = 14'h12D8;
            14'd13913: out = 14'h12D7;
            14'd13914: out = 14'h12D7;
            14'd13915: out = 14'h12D7;
            14'd13916: out = 14'h12D6;
            14'd13917: out = 14'h12D6;
            14'd13918: out = 14'h12D6;
            14'd13919: out = 14'h12D5;
            14'd13920: out = 14'h12D5;
            14'd13921: out = 14'h12D5;
            14'd13922: out = 14'h12D4;
            14'd13923: out = 14'h12D4;
            14'd13924: out = 14'h12D4;
            14'd13925: out = 14'h12D3;
            14'd13926: out = 14'h12D3;
            14'd13927: out = 14'h12D3;
            14'd13928: out = 14'h12D2;
            14'd13929: out = 14'h12D2;
            14'd13930: out = 14'h12D2;
            14'd13931: out = 14'h12D1;
            14'd13932: out = 14'h12D1;
            14'd13933: out = 14'h12D1;
            14'd13934: out = 14'h12D0;
            14'd13935: out = 14'h12D0;
            14'd13936: out = 14'h12D0;
            14'd13937: out = 14'h12CF;
            14'd13938: out = 14'h12CF;
            14'd13939: out = 14'h12CE;
            14'd13940: out = 14'h12CE;
            14'd13941: out = 14'h12CE;
            14'd13942: out = 14'h12CD;
            14'd13943: out = 14'h12CD;
            14'd13944: out = 14'h12CD;
            14'd13945: out = 14'h12CC;
            14'd13946: out = 14'h12CC;
            14'd13947: out = 14'h12CC;
            14'd13948: out = 14'h12CB;
            14'd13949: out = 14'h12CB;
            14'd13950: out = 14'h12CB;
            14'd13951: out = 14'h12CA;
            14'd13952: out = 14'h12CA;
            14'd13953: out = 14'h12CA;
            14'd13954: out = 14'h12C9;
            14'd13955: out = 14'h12C9;
            14'd13956: out = 14'h12C9;
            14'd13957: out = 14'h12C8;
            14'd13958: out = 14'h12C8;
            14'd13959: out = 14'h12C8;
            14'd13960: out = 14'h12C7;
            14'd13961: out = 14'h12C7;
            14'd13962: out = 14'h12C7;
            14'd13963: out = 14'h12C6;
            14'd13964: out = 14'h12C6;
            14'd13965: out = 14'h12C6;
            14'd13966: out = 14'h12C5;
            14'd13967: out = 14'h12C5;
            14'd13968: out = 14'h12C4;
            14'd13969: out = 14'h12C4;
            14'd13970: out = 14'h12C4;
            14'd13971: out = 14'h12C3;
            14'd13972: out = 14'h12C3;
            14'd13973: out = 14'h12C3;
            14'd13974: out = 14'h12C2;
            14'd13975: out = 14'h12C2;
            14'd13976: out = 14'h12C2;
            14'd13977: out = 14'h12C1;
            14'd13978: out = 14'h12C1;
            14'd13979: out = 14'h12C1;
            14'd13980: out = 14'h12C0;
            14'd13981: out = 14'h12C0;
            14'd13982: out = 14'h12C0;
            14'd13983: out = 14'h12BF;
            14'd13984: out = 14'h12BF;
            14'd13985: out = 14'h12BF;
            14'd13986: out = 14'h12BE;
            14'd13987: out = 14'h12BE;
            14'd13988: out = 14'h12BE;
            14'd13989: out = 14'h12BD;
            14'd13990: out = 14'h12BD;
            14'd13991: out = 14'h12BD;
            14'd13992: out = 14'h12BC;
            14'd13993: out = 14'h12BC;
            14'd13994: out = 14'h12BC;
            14'd13995: out = 14'h12BB;
            14'd13996: out = 14'h12BB;
            14'd13997: out = 14'h12BB;
            14'd13998: out = 14'h12BA;
            14'd13999: out = 14'h12BA;
            14'd14000: out = 14'h12B9;
            14'd14001: out = 14'h12B9;
            14'd14002: out = 14'h12B9;
            14'd14003: out = 14'h12B8;
            14'd14004: out = 14'h12B8;
            14'd14005: out = 14'h12B8;
            14'd14006: out = 14'h12B7;
            14'd14007: out = 14'h12B7;
            14'd14008: out = 14'h12B7;
            14'd14009: out = 14'h12B6;
            14'd14010: out = 14'h12B6;
            14'd14011: out = 14'h12B6;
            14'd14012: out = 14'h12B5;
            14'd14013: out = 14'h12B5;
            14'd14014: out = 14'h12B5;
            14'd14015: out = 14'h12B4;
            14'd14016: out = 14'h12B4;
            14'd14017: out = 14'h12B4;
            14'd14018: out = 14'h12B3;
            14'd14019: out = 14'h12B3;
            14'd14020: out = 14'h12B3;
            14'd14021: out = 14'h12B2;
            14'd14022: out = 14'h12B2;
            14'd14023: out = 14'h12B2;
            14'd14024: out = 14'h12B1;
            14'd14025: out = 14'h12B1;
            14'd14026: out = 14'h12B1;
            14'd14027: out = 14'h12B0;
            14'd14028: out = 14'h12B0;
            14'd14029: out = 14'h12B0;
            14'd14030: out = 14'h12AF;
            14'd14031: out = 14'h12AF;
            14'd14032: out = 14'h12AF;
            14'd14033: out = 14'h12AE;
            14'd14034: out = 14'h12AE;
            14'd14035: out = 14'h12AE;
            14'd14036: out = 14'h12AD;
            14'd14037: out = 14'h12AD;
            14'd14038: out = 14'h12AD;
            14'd14039: out = 14'h12AC;
            14'd14040: out = 14'h12AC;
            14'd14041: out = 14'h12AB;
            14'd14042: out = 14'h12AB;
            14'd14043: out = 14'h12AB;
            14'd14044: out = 14'h12AA;
            14'd14045: out = 14'h12AA;
            14'd14046: out = 14'h12AA;
            14'd14047: out = 14'h12A9;
            14'd14048: out = 14'h12A9;
            14'd14049: out = 14'h12A9;
            14'd14050: out = 14'h12A8;
            14'd14051: out = 14'h12A8;
            14'd14052: out = 14'h12A8;
            14'd14053: out = 14'h12A7;
            14'd14054: out = 14'h12A7;
            14'd14055: out = 14'h12A7;
            14'd14056: out = 14'h12A6;
            14'd14057: out = 14'h12A6;
            14'd14058: out = 14'h12A6;
            14'd14059: out = 14'h12A5;
            14'd14060: out = 14'h12A5;
            14'd14061: out = 14'h12A5;
            14'd14062: out = 14'h12A4;
            14'd14063: out = 14'h12A4;
            14'd14064: out = 14'h12A4;
            14'd14065: out = 14'h12A3;
            14'd14066: out = 14'h12A3;
            14'd14067: out = 14'h12A3;
            14'd14068: out = 14'h12A2;
            14'd14069: out = 14'h12A2;
            14'd14070: out = 14'h12A2;
            14'd14071: out = 14'h12A1;
            14'd14072: out = 14'h12A1;
            14'd14073: out = 14'h12A1;
            14'd14074: out = 14'h12A0;
            14'd14075: out = 14'h12A0;
            14'd14076: out = 14'h12A0;
            14'd14077: out = 14'h129F;
            14'd14078: out = 14'h129F;
            14'd14079: out = 14'h129F;
            14'd14080: out = 14'h129E;
            14'd14081: out = 14'h129E;
            14'd14082: out = 14'h129E;
            14'd14083: out = 14'h129D;
            14'd14084: out = 14'h129D;
            14'd14085: out = 14'h129D;
            14'd14086: out = 14'h129C;
            14'd14087: out = 14'h129C;
            14'd14088: out = 14'h129C;
            14'd14089: out = 14'h129B;
            14'd14090: out = 14'h129B;
            14'd14091: out = 14'h129B;
            14'd14092: out = 14'h129A;
            14'd14093: out = 14'h129A;
            14'd14094: out = 14'h129A;
            14'd14095: out = 14'h1299;
            14'd14096: out = 14'h1299;
            14'd14097: out = 14'h1299;
            14'd14098: out = 14'h1298;
            14'd14099: out = 14'h1298;
            14'd14100: out = 14'h1297;
            14'd14101: out = 14'h1297;
            14'd14102: out = 14'h1297;
            14'd14103: out = 14'h1296;
            14'd14104: out = 14'h1296;
            14'd14105: out = 14'h1296;
            14'd14106: out = 14'h1295;
            14'd14107: out = 14'h1295;
            14'd14108: out = 14'h1295;
            14'd14109: out = 14'h1294;
            14'd14110: out = 14'h1294;
            14'd14111: out = 14'h1294;
            14'd14112: out = 14'h1293;
            14'd14113: out = 14'h1293;
            14'd14114: out = 14'h1293;
            14'd14115: out = 14'h1292;
            14'd14116: out = 14'h1292;
            14'd14117: out = 14'h1292;
            14'd14118: out = 14'h1291;
            14'd14119: out = 14'h1291;
            14'd14120: out = 14'h1291;
            14'd14121: out = 14'h1290;
            14'd14122: out = 14'h1290;
            14'd14123: out = 14'h1290;
            14'd14124: out = 14'h128F;
            14'd14125: out = 14'h128F;
            14'd14126: out = 14'h128F;
            14'd14127: out = 14'h128E;
            14'd14128: out = 14'h128E;
            14'd14129: out = 14'h128E;
            14'd14130: out = 14'h128D;
            14'd14131: out = 14'h128D;
            14'd14132: out = 14'h128D;
            14'd14133: out = 14'h128C;
            14'd14134: out = 14'h128C;
            14'd14135: out = 14'h128C;
            14'd14136: out = 14'h128B;
            14'd14137: out = 14'h128B;
            14'd14138: out = 14'h128B;
            14'd14139: out = 14'h128A;
            14'd14140: out = 14'h128A;
            14'd14141: out = 14'h128A;
            14'd14142: out = 14'h1289;
            14'd14143: out = 14'h1289;
            14'd14144: out = 14'h1289;
            14'd14145: out = 14'h1288;
            14'd14146: out = 14'h1288;
            14'd14147: out = 14'h1288;
            14'd14148: out = 14'h1287;
            14'd14149: out = 14'h1287;
            14'd14150: out = 14'h1287;
            14'd14151: out = 14'h1286;
            14'd14152: out = 14'h1286;
            14'd14153: out = 14'h1286;
            14'd14154: out = 14'h1285;
            14'd14155: out = 14'h1285;
            14'd14156: out = 14'h1285;
            14'd14157: out = 14'h1284;
            14'd14158: out = 14'h1284;
            14'd14159: out = 14'h1284;
            14'd14160: out = 14'h1283;
            14'd14161: out = 14'h1283;
            14'd14162: out = 14'h1283;
            14'd14163: out = 14'h1282;
            14'd14164: out = 14'h1282;
            14'd14165: out = 14'h1282;
            14'd14166: out = 14'h1281;
            14'd14167: out = 14'h1281;
            14'd14168: out = 14'h1281;
            14'd14169: out = 14'h1280;
            14'd14170: out = 14'h1280;
            14'd14171: out = 14'h1280;
            14'd14172: out = 14'h127F;
            14'd14173: out = 14'h127F;
            14'd14174: out = 14'h127F;
            14'd14175: out = 14'h127E;
            14'd14176: out = 14'h127E;
            14'd14177: out = 14'h127E;
            14'd14178: out = 14'h127D;
            14'd14179: out = 14'h127D;
            14'd14180: out = 14'h127D;
            14'd14181: out = 14'h127C;
            14'd14182: out = 14'h127C;
            14'd14183: out = 14'h127C;
            14'd14184: out = 14'h127B;
            14'd14185: out = 14'h127B;
            14'd14186: out = 14'h127B;
            14'd14187: out = 14'h127A;
            14'd14188: out = 14'h127A;
            14'd14189: out = 14'h127A;
            14'd14190: out = 14'h1279;
            14'd14191: out = 14'h1279;
            14'd14192: out = 14'h1279;
            14'd14193: out = 14'h1278;
            14'd14194: out = 14'h1278;
            14'd14195: out = 14'h1278;
            14'd14196: out = 14'h1277;
            14'd14197: out = 14'h1277;
            14'd14198: out = 14'h1277;
            14'd14199: out = 14'h1276;
            14'd14200: out = 14'h1276;
            14'd14201: out = 14'h1276;
            14'd14202: out = 14'h1275;
            14'd14203: out = 14'h1275;
            14'd14204: out = 14'h1275;
            14'd14205: out = 14'h1274;
            14'd14206: out = 14'h1274;
            14'd14207: out = 14'h1274;
            14'd14208: out = 14'h1273;
            14'd14209: out = 14'h1273;
            14'd14210: out = 14'h1273;
            14'd14211: out = 14'h1272;
            14'd14212: out = 14'h1272;
            14'd14213: out = 14'h1272;
            14'd14214: out = 14'h1271;
            14'd14215: out = 14'h1271;
            14'd14216: out = 14'h1271;
            14'd14217: out = 14'h1270;
            14'd14218: out = 14'h1270;
            14'd14219: out = 14'h1270;
            14'd14220: out = 14'h126F;
            14'd14221: out = 14'h126F;
            14'd14222: out = 14'h126F;
            14'd14223: out = 14'h126E;
            14'd14224: out = 14'h126E;
            14'd14225: out = 14'h126E;
            14'd14226: out = 14'h126D;
            14'd14227: out = 14'h126D;
            14'd14228: out = 14'h126D;
            14'd14229: out = 14'h126C;
            14'd14230: out = 14'h126C;
            14'd14231: out = 14'h126C;
            14'd14232: out = 14'h126B;
            14'd14233: out = 14'h126B;
            14'd14234: out = 14'h126B;
            14'd14235: out = 14'h126A;
            14'd14236: out = 14'h126A;
            14'd14237: out = 14'h126A;
            14'd14238: out = 14'h1269;
            14'd14239: out = 14'h1269;
            14'd14240: out = 14'h1269;
            14'd14241: out = 14'h1268;
            14'd14242: out = 14'h1268;
            14'd14243: out = 14'h1268;
            14'd14244: out = 14'h1267;
            14'd14245: out = 14'h1267;
            14'd14246: out = 14'h1267;
            14'd14247: out = 14'h1266;
            14'd14248: out = 14'h1266;
            14'd14249: out = 14'h1266;
            14'd14250: out = 14'h1265;
            14'd14251: out = 14'h1265;
            14'd14252: out = 14'h1265;
            14'd14253: out = 14'h1264;
            14'd14254: out = 14'h1264;
            14'd14255: out = 14'h1264;
            14'd14256: out = 14'h1263;
            14'd14257: out = 14'h1263;
            14'd14258: out = 14'h1263;
            14'd14259: out = 14'h1262;
            14'd14260: out = 14'h1262;
            14'd14261: out = 14'h1262;
            14'd14262: out = 14'h1261;
            14'd14263: out = 14'h1261;
            14'd14264: out = 14'h1261;
            14'd14265: out = 14'h1260;
            14'd14266: out = 14'h1260;
            14'd14267: out = 14'h1260;
            14'd14268: out = 14'h125F;
            14'd14269: out = 14'h125F;
            14'd14270: out = 14'h125F;
            14'd14271: out = 14'h125E;
            14'd14272: out = 14'h125E;
            14'd14273: out = 14'h125E;
            14'd14274: out = 14'h125D;
            14'd14275: out = 14'h125D;
            14'd14276: out = 14'h125D;
            14'd14277: out = 14'h125C;
            14'd14278: out = 14'h125C;
            14'd14279: out = 14'h125C;
            14'd14280: out = 14'h125C;
            14'd14281: out = 14'h125B;
            14'd14282: out = 14'h125B;
            14'd14283: out = 14'h125B;
            14'd14284: out = 14'h125A;
            14'd14285: out = 14'h125A;
            14'd14286: out = 14'h125A;
            14'd14287: out = 14'h1259;
            14'd14288: out = 14'h1259;
            14'd14289: out = 14'h1259;
            14'd14290: out = 14'h1258;
            14'd14291: out = 14'h1258;
            14'd14292: out = 14'h1258;
            14'd14293: out = 14'h1257;
            14'd14294: out = 14'h1257;
            14'd14295: out = 14'h1257;
            14'd14296: out = 14'h1256;
            14'd14297: out = 14'h1256;
            14'd14298: out = 14'h1256;
            14'd14299: out = 14'h1255;
            14'd14300: out = 14'h1255;
            14'd14301: out = 14'h1255;
            14'd14302: out = 14'h1254;
            14'd14303: out = 14'h1254;
            14'd14304: out = 14'h1254;
            14'd14305: out = 14'h1253;
            14'd14306: out = 14'h1253;
            14'd14307: out = 14'h1253;
            14'd14308: out = 14'h1252;
            14'd14309: out = 14'h1252;
            14'd14310: out = 14'h1252;
            14'd14311: out = 14'h1251;
            14'd14312: out = 14'h1251;
            14'd14313: out = 14'h1251;
            14'd14314: out = 14'h1250;
            14'd14315: out = 14'h1250;
            14'd14316: out = 14'h1250;
            14'd14317: out = 14'h124F;
            14'd14318: out = 14'h124F;
            14'd14319: out = 14'h124F;
            14'd14320: out = 14'h124E;
            14'd14321: out = 14'h124E;
            14'd14322: out = 14'h124E;
            14'd14323: out = 14'h124D;
            14'd14324: out = 14'h124D;
            14'd14325: out = 14'h124D;
            14'd14326: out = 14'h124C;
            14'd14327: out = 14'h124C;
            14'd14328: out = 14'h124C;
            14'd14329: out = 14'h124B;
            14'd14330: out = 14'h124B;
            14'd14331: out = 14'h124B;
            14'd14332: out = 14'h124A;
            14'd14333: out = 14'h124A;
            14'd14334: out = 14'h124A;
            14'd14335: out = 14'h1249;
            14'd14336: out = 14'h1249;
            14'd14337: out = 14'h1249;
            14'd14338: out = 14'h1248;
            14'd14339: out = 14'h1248;
            14'd14340: out = 14'h1248;
            14'd14341: out = 14'h1248;
            14'd14342: out = 14'h1247;
            14'd14343: out = 14'h1247;
            14'd14344: out = 14'h1247;
            14'd14345: out = 14'h1246;
            14'd14346: out = 14'h1246;
            14'd14347: out = 14'h1246;
            14'd14348: out = 14'h1245;
            14'd14349: out = 14'h1245;
            14'd14350: out = 14'h1245;
            14'd14351: out = 14'h1244;
            14'd14352: out = 14'h1244;
            14'd14353: out = 14'h1244;
            14'd14354: out = 14'h1243;
            14'd14355: out = 14'h1243;
            14'd14356: out = 14'h1243;
            14'd14357: out = 14'h1242;
            14'd14358: out = 14'h1242;
            14'd14359: out = 14'h1242;
            14'd14360: out = 14'h1241;
            14'd14361: out = 14'h1241;
            14'd14362: out = 14'h1241;
            14'd14363: out = 14'h1240;
            14'd14364: out = 14'h1240;
            14'd14365: out = 14'h1240;
            14'd14366: out = 14'h123F;
            14'd14367: out = 14'h123F;
            14'd14368: out = 14'h123F;
            14'd14369: out = 14'h123E;
            14'd14370: out = 14'h123E;
            14'd14371: out = 14'h123E;
            14'd14372: out = 14'h123D;
            14'd14373: out = 14'h123D;
            14'd14374: out = 14'h123D;
            14'd14375: out = 14'h123C;
            14'd14376: out = 14'h123C;
            14'd14377: out = 14'h123C;
            14'd14378: out = 14'h123B;
            14'd14379: out = 14'h123B;
            14'd14380: out = 14'h123B;
            14'd14381: out = 14'h123A;
            14'd14382: out = 14'h123A;
            14'd14383: out = 14'h123A;
            14'd14384: out = 14'h123A;
            14'd14385: out = 14'h1239;
            14'd14386: out = 14'h1239;
            14'd14387: out = 14'h1239;
            14'd14388: out = 14'h1238;
            14'd14389: out = 14'h1238;
            14'd14390: out = 14'h1238;
            14'd14391: out = 14'h1237;
            14'd14392: out = 14'h1237;
            14'd14393: out = 14'h1237;
            14'd14394: out = 14'h1236;
            14'd14395: out = 14'h1236;
            14'd14396: out = 14'h1236;
            14'd14397: out = 14'h1235;
            14'd14398: out = 14'h1235;
            14'd14399: out = 14'h1235;
            14'd14400: out = 14'h1234;
            14'd14401: out = 14'h1234;
            14'd14402: out = 14'h1234;
            14'd14403: out = 14'h1233;
            14'd14404: out = 14'h1233;
            14'd14405: out = 14'h1233;
            14'd14406: out = 14'h1232;
            14'd14407: out = 14'h1232;
            14'd14408: out = 14'h1232;
            14'd14409: out = 14'h1231;
            14'd14410: out = 14'h1231;
            14'd14411: out = 14'h1231;
            14'd14412: out = 14'h1230;
            14'd14413: out = 14'h1230;
            14'd14414: out = 14'h1230;
            14'd14415: out = 14'h122F;
            14'd14416: out = 14'h122F;
            14'd14417: out = 14'h122F;
            14'd14418: out = 14'h122F;
            14'd14419: out = 14'h122E;
            14'd14420: out = 14'h122E;
            14'd14421: out = 14'h122E;
            14'd14422: out = 14'h122D;
            14'd14423: out = 14'h122D;
            14'd14424: out = 14'h122D;
            14'd14425: out = 14'h122C;
            14'd14426: out = 14'h122C;
            14'd14427: out = 14'h122C;
            14'd14428: out = 14'h122B;
            14'd14429: out = 14'h122B;
            14'd14430: out = 14'h122B;
            14'd14431: out = 14'h122A;
            14'd14432: out = 14'h122A;
            14'd14433: out = 14'h122A;
            14'd14434: out = 14'h1229;
            14'd14435: out = 14'h1229;
            14'd14436: out = 14'h1229;
            14'd14437: out = 14'h1228;
            14'd14438: out = 14'h1228;
            14'd14439: out = 14'h1228;
            14'd14440: out = 14'h1227;
            14'd14441: out = 14'h1227;
            14'd14442: out = 14'h1227;
            14'd14443: out = 14'h1226;
            14'd14444: out = 14'h1226;
            14'd14445: out = 14'h1226;
            14'd14446: out = 14'h1225;
            14'd14447: out = 14'h1225;
            14'd14448: out = 14'h1225;
            14'd14449: out = 14'h1225;
            14'd14450: out = 14'h1224;
            14'd14451: out = 14'h1224;
            14'd14452: out = 14'h1224;
            14'd14453: out = 14'h1223;
            14'd14454: out = 14'h1223;
            14'd14455: out = 14'h1223;
            14'd14456: out = 14'h1222;
            14'd14457: out = 14'h1222;
            14'd14458: out = 14'h1222;
            14'd14459: out = 14'h1221;
            14'd14460: out = 14'h1221;
            14'd14461: out = 14'h1221;
            14'd14462: out = 14'h1220;
            14'd14463: out = 14'h1220;
            14'd14464: out = 14'h1220;
            14'd14465: out = 14'h121F;
            14'd14466: out = 14'h121F;
            14'd14467: out = 14'h121F;
            14'd14468: out = 14'h121E;
            14'd14469: out = 14'h121E;
            14'd14470: out = 14'h121E;
            14'd14471: out = 14'h121D;
            14'd14472: out = 14'h121D;
            14'd14473: out = 14'h121D;
            14'd14474: out = 14'h121D;
            14'd14475: out = 14'h121C;
            14'd14476: out = 14'h121C;
            14'd14477: out = 14'h121C;
            14'd14478: out = 14'h121B;
            14'd14479: out = 14'h121B;
            14'd14480: out = 14'h121B;
            14'd14481: out = 14'h121A;
            14'd14482: out = 14'h121A;
            14'd14483: out = 14'h121A;
            14'd14484: out = 14'h1219;
            14'd14485: out = 14'h1219;
            14'd14486: out = 14'h1219;
            14'd14487: out = 14'h1218;
            14'd14488: out = 14'h1218;
            14'd14489: out = 14'h1218;
            14'd14490: out = 14'h1217;
            14'd14491: out = 14'h1217;
            14'd14492: out = 14'h1217;
            14'd14493: out = 14'h1216;
            14'd14494: out = 14'h1216;
            14'd14495: out = 14'h1216;
            14'd14496: out = 14'h1215;
            14'd14497: out = 14'h1215;
            14'd14498: out = 14'h1215;
            14'd14499: out = 14'h1215;
            14'd14500: out = 14'h1214;
            14'd14501: out = 14'h1214;
            14'd14502: out = 14'h1214;
            14'd14503: out = 14'h1213;
            14'd14504: out = 14'h1213;
            14'd14505: out = 14'h1213;
            14'd14506: out = 14'h1212;
            14'd14507: out = 14'h1212;
            14'd14508: out = 14'h1212;
            14'd14509: out = 14'h1211;
            14'd14510: out = 14'h1211;
            14'd14511: out = 14'h1211;
            14'd14512: out = 14'h1210;
            14'd14513: out = 14'h1210;
            14'd14514: out = 14'h1210;
            14'd14515: out = 14'h120F;
            14'd14516: out = 14'h120F;
            14'd14517: out = 14'h120F;
            14'd14518: out = 14'h120E;
            14'd14519: out = 14'h120E;
            14'd14520: out = 14'h120E;
            14'd14521: out = 14'h120E;
            14'd14522: out = 14'h120D;
            14'd14523: out = 14'h120D;
            14'd14524: out = 14'h120D;
            14'd14525: out = 14'h120C;
            14'd14526: out = 14'h120C;
            14'd14527: out = 14'h120C;
            14'd14528: out = 14'h120B;
            14'd14529: out = 14'h120B;
            14'd14530: out = 14'h120B;
            14'd14531: out = 14'h120A;
            14'd14532: out = 14'h120A;
            14'd14533: out = 14'h120A;
            14'd14534: out = 14'h1209;
            14'd14535: out = 14'h1209;
            14'd14536: out = 14'h1209;
            14'd14537: out = 14'h1208;
            14'd14538: out = 14'h1208;
            14'd14539: out = 14'h1208;
            14'd14540: out = 14'h1207;
            14'd14541: out = 14'h1207;
            14'd14542: out = 14'h1207;
            14'd14543: out = 14'h1207;
            14'd14544: out = 14'h1206;
            14'd14545: out = 14'h1206;
            14'd14546: out = 14'h1206;
            14'd14547: out = 14'h1205;
            14'd14548: out = 14'h1205;
            14'd14549: out = 14'h1205;
            14'd14550: out = 14'h1204;
            14'd14551: out = 14'h1204;
            14'd14552: out = 14'h1204;
            14'd14553: out = 14'h1203;
            14'd14554: out = 14'h1203;
            14'd14555: out = 14'h1203;
            14'd14556: out = 14'h1202;
            14'd14557: out = 14'h1202;
            14'd14558: out = 14'h1202;
            14'd14559: out = 14'h1201;
            14'd14560: out = 14'h1201;
            14'd14561: out = 14'h1201;
            14'd14562: out = 14'h1200;
            14'd14563: out = 14'h1200;
            14'd14564: out = 14'h1200;
            14'd14565: out = 14'h1200;
            14'd14566: out = 14'h11FF;
            14'd14567: out = 14'h11FF;
            14'd14568: out = 14'h11FF;
            14'd14569: out = 14'h11FE;
            14'd14570: out = 14'h11FE;
            14'd14571: out = 14'h11FE;
            14'd14572: out = 14'h11FD;
            14'd14573: out = 14'h11FD;
            14'd14574: out = 14'h11FD;
            14'd14575: out = 14'h11FC;
            14'd14576: out = 14'h11FC;
            14'd14577: out = 14'h11FC;
            14'd14578: out = 14'h11FB;
            14'd14579: out = 14'h11FB;
            14'd14580: out = 14'h11FB;
            14'd14581: out = 14'h11FA;
            14'd14582: out = 14'h11FA;
            14'd14583: out = 14'h11FA;
            14'd14584: out = 14'h11FA;
            14'd14585: out = 14'h11F9;
            14'd14586: out = 14'h11F9;
            14'd14587: out = 14'h11F9;
            14'd14588: out = 14'h11F8;
            14'd14589: out = 14'h11F8;
            14'd14590: out = 14'h11F8;
            14'd14591: out = 14'h11F7;
            14'd14592: out = 14'h11F7;
            14'd14593: out = 14'h11F7;
            14'd14594: out = 14'h11F6;
            14'd14595: out = 14'h11F6;
            14'd14596: out = 14'h11F6;
            14'd14597: out = 14'h11F5;
            14'd14598: out = 14'h11F5;
            14'd14599: out = 14'h11F5;
            14'd14600: out = 14'h11F4;
            14'd14601: out = 14'h11F4;
            14'd14602: out = 14'h11F4;
            14'd14603: out = 14'h11F4;
            14'd14604: out = 14'h11F3;
            14'd14605: out = 14'h11F3;
            14'd14606: out = 14'h11F3;
            14'd14607: out = 14'h11F2;
            14'd14608: out = 14'h11F2;
            14'd14609: out = 14'h11F2;
            14'd14610: out = 14'h11F1;
            14'd14611: out = 14'h11F1;
            14'd14612: out = 14'h11F1;
            14'd14613: out = 14'h11F0;
            14'd14614: out = 14'h11F0;
            14'd14615: out = 14'h11F0;
            14'd14616: out = 14'h11EF;
            14'd14617: out = 14'h11EF;
            14'd14618: out = 14'h11EF;
            14'd14619: out = 14'h11EF;
            14'd14620: out = 14'h11EE;
            14'd14621: out = 14'h11EE;
            14'd14622: out = 14'h11EE;
            14'd14623: out = 14'h11ED;
            14'd14624: out = 14'h11ED;
            14'd14625: out = 14'h11ED;
            14'd14626: out = 14'h11EC;
            14'd14627: out = 14'h11EC;
            14'd14628: out = 14'h11EC;
            14'd14629: out = 14'h11EB;
            14'd14630: out = 14'h11EB;
            14'd14631: out = 14'h11EB;
            14'd14632: out = 14'h11EA;
            14'd14633: out = 14'h11EA;
            14'd14634: out = 14'h11EA;
            14'd14635: out = 14'h11EA;
            14'd14636: out = 14'h11E9;
            14'd14637: out = 14'h11E9;
            14'd14638: out = 14'h11E9;
            14'd14639: out = 14'h11E8;
            14'd14640: out = 14'h11E8;
            14'd14641: out = 14'h11E8;
            14'd14642: out = 14'h11E7;
            14'd14643: out = 14'h11E7;
            14'd14644: out = 14'h11E7;
            14'd14645: out = 14'h11E6;
            14'd14646: out = 14'h11E6;
            14'd14647: out = 14'h11E6;
            14'd14648: out = 14'h11E5;
            14'd14649: out = 14'h11E5;
            14'd14650: out = 14'h11E5;
            14'd14651: out = 14'h11E4;
            14'd14652: out = 14'h11E4;
            14'd14653: out = 14'h11E4;
            14'd14654: out = 14'h11E4;
            14'd14655: out = 14'h11E3;
            14'd14656: out = 14'h11E3;
            14'd14657: out = 14'h11E3;
            14'd14658: out = 14'h11E2;
            14'd14659: out = 14'h11E2;
            14'd14660: out = 14'h11E2;
            14'd14661: out = 14'h11E1;
            14'd14662: out = 14'h11E1;
            14'd14663: out = 14'h11E1;
            14'd14664: out = 14'h11E0;
            14'd14665: out = 14'h11E0;
            14'd14666: out = 14'h11E0;
            14'd14667: out = 14'h11E0;
            14'd14668: out = 14'h11DF;
            14'd14669: out = 14'h11DF;
            14'd14670: out = 14'h11DF;
            14'd14671: out = 14'h11DE;
            14'd14672: out = 14'h11DE;
            14'd14673: out = 14'h11DE;
            14'd14674: out = 14'h11DD;
            14'd14675: out = 14'h11DD;
            14'd14676: out = 14'h11DD;
            14'd14677: out = 14'h11DC;
            14'd14678: out = 14'h11DC;
            14'd14679: out = 14'h11DC;
            14'd14680: out = 14'h11DB;
            14'd14681: out = 14'h11DB;
            14'd14682: out = 14'h11DB;
            14'd14683: out = 14'h11DB;
            14'd14684: out = 14'h11DA;
            14'd14685: out = 14'h11DA;
            14'd14686: out = 14'h11DA;
            14'd14687: out = 14'h11D9;
            14'd14688: out = 14'h11D9;
            14'd14689: out = 14'h11D9;
            14'd14690: out = 14'h11D8;
            14'd14691: out = 14'h11D8;
            14'd14692: out = 14'h11D8;
            14'd14693: out = 14'h11D7;
            14'd14694: out = 14'h11D7;
            14'd14695: out = 14'h11D7;
            14'd14696: out = 14'h11D6;
            14'd14697: out = 14'h11D6;
            14'd14698: out = 14'h11D6;
            14'd14699: out = 14'h11D6;
            14'd14700: out = 14'h11D5;
            14'd14701: out = 14'h11D5;
            14'd14702: out = 14'h11D5;
            14'd14703: out = 14'h11D4;
            14'd14704: out = 14'h11D4;
            14'd14705: out = 14'h11D4;
            14'd14706: out = 14'h11D3;
            14'd14707: out = 14'h11D3;
            14'd14708: out = 14'h11D3;
            14'd14709: out = 14'h11D2;
            14'd14710: out = 14'h11D2;
            14'd14711: out = 14'h11D2;
            14'd14712: out = 14'h11D2;
            14'd14713: out = 14'h11D1;
            14'd14714: out = 14'h11D1;
            14'd14715: out = 14'h11D1;
            14'd14716: out = 14'h11D0;
            14'd14717: out = 14'h11D0;
            14'd14718: out = 14'h11D0;
            14'd14719: out = 14'h11CF;
            14'd14720: out = 14'h11CF;
            14'd14721: out = 14'h11CF;
            14'd14722: out = 14'h11CE;
            14'd14723: out = 14'h11CE;
            14'd14724: out = 14'h11CE;
            14'd14725: out = 14'h11CD;
            14'd14726: out = 14'h11CD;
            14'd14727: out = 14'h11CD;
            14'd14728: out = 14'h11CD;
            14'd14729: out = 14'h11CC;
            14'd14730: out = 14'h11CC;
            14'd14731: out = 14'h11CC;
            14'd14732: out = 14'h11CB;
            14'd14733: out = 14'h11CB;
            14'd14734: out = 14'h11CB;
            14'd14735: out = 14'h11CA;
            14'd14736: out = 14'h11CA;
            14'd14737: out = 14'h11CA;
            14'd14738: out = 14'h11C9;
            14'd14739: out = 14'h11C9;
            14'd14740: out = 14'h11C9;
            14'd14741: out = 14'h11C9;
            14'd14742: out = 14'h11C8;
            14'd14743: out = 14'h11C8;
            14'd14744: out = 14'h11C8;
            14'd14745: out = 14'h11C7;
            14'd14746: out = 14'h11C7;
            14'd14747: out = 14'h11C7;
            14'd14748: out = 14'h11C6;
            14'd14749: out = 14'h11C6;
            14'd14750: out = 14'h11C6;
            14'd14751: out = 14'h11C5;
            14'd14752: out = 14'h11C5;
            14'd14753: out = 14'h11C5;
            14'd14754: out = 14'h11C5;
            14'd14755: out = 14'h11C4;
            14'd14756: out = 14'h11C4;
            14'd14757: out = 14'h11C4;
            14'd14758: out = 14'h11C3;
            14'd14759: out = 14'h11C3;
            14'd14760: out = 14'h11C3;
            14'd14761: out = 14'h11C2;
            14'd14762: out = 14'h11C2;
            14'd14763: out = 14'h11C2;
            14'd14764: out = 14'h11C1;
            14'd14765: out = 14'h11C1;
            14'd14766: out = 14'h11C1;
            14'd14767: out = 14'h11C1;
            14'd14768: out = 14'h11C0;
            14'd14769: out = 14'h11C0;
            14'd14770: out = 14'h11C0;
            14'd14771: out = 14'h11BF;
            14'd14772: out = 14'h11BF;
            14'd14773: out = 14'h11BF;
            14'd14774: out = 14'h11BE;
            14'd14775: out = 14'h11BE;
            14'd14776: out = 14'h11BE;
            14'd14777: out = 14'h11BD;
            14'd14778: out = 14'h11BD;
            14'd14779: out = 14'h11BD;
            14'd14780: out = 14'h11BD;
            14'd14781: out = 14'h11BC;
            14'd14782: out = 14'h11BC;
            14'd14783: out = 14'h11BC;
            14'd14784: out = 14'h11BB;
            14'd14785: out = 14'h11BB;
            14'd14786: out = 14'h11BB;
            14'd14787: out = 14'h11BA;
            14'd14788: out = 14'h11BA;
            14'd14789: out = 14'h11BA;
            14'd14790: out = 14'h11B9;
            14'd14791: out = 14'h11B9;
            14'd14792: out = 14'h11B9;
            14'd14793: out = 14'h11B9;
            14'd14794: out = 14'h11B8;
            14'd14795: out = 14'h11B8;
            14'd14796: out = 14'h11B8;
            14'd14797: out = 14'h11B7;
            14'd14798: out = 14'h11B7;
            14'd14799: out = 14'h11B7;
            14'd14800: out = 14'h11B6;
            14'd14801: out = 14'h11B6;
            14'd14802: out = 14'h11B6;
            14'd14803: out = 14'h11B5;
            14'd14804: out = 14'h11B5;
            14'd14805: out = 14'h11B5;
            14'd14806: out = 14'h11B5;
            14'd14807: out = 14'h11B4;
            14'd14808: out = 14'h11B4;
            14'd14809: out = 14'h11B4;
            14'd14810: out = 14'h11B3;
            14'd14811: out = 14'h11B3;
            14'd14812: out = 14'h11B3;
            14'd14813: out = 14'h11B2;
            14'd14814: out = 14'h11B2;
            14'd14815: out = 14'h11B2;
            14'd14816: out = 14'h11B1;
            14'd14817: out = 14'h11B1;
            14'd14818: out = 14'h11B1;
            14'd14819: out = 14'h11B1;
            14'd14820: out = 14'h11B0;
            14'd14821: out = 14'h11B0;
            14'd14822: out = 14'h11B0;
            14'd14823: out = 14'h11AF;
            14'd14824: out = 14'h11AF;
            14'd14825: out = 14'h11AF;
            14'd14826: out = 14'h11AE;
            14'd14827: out = 14'h11AE;
            14'd14828: out = 14'h11AE;
            14'd14829: out = 14'h11AE;
            14'd14830: out = 14'h11AD;
            14'd14831: out = 14'h11AD;
            14'd14832: out = 14'h11AD;
            14'd14833: out = 14'h11AC;
            14'd14834: out = 14'h11AC;
            14'd14835: out = 14'h11AC;
            14'd14836: out = 14'h11AB;
            14'd14837: out = 14'h11AB;
            14'd14838: out = 14'h11AB;
            14'd14839: out = 14'h11AA;
            14'd14840: out = 14'h11AA;
            14'd14841: out = 14'h11AA;
            14'd14842: out = 14'h11AA;
            14'd14843: out = 14'h11A9;
            14'd14844: out = 14'h11A9;
            14'd14845: out = 14'h11A9;
            14'd14846: out = 14'h11A8;
            14'd14847: out = 14'h11A8;
            14'd14848: out = 14'h11A8;
            14'd14849: out = 14'h11A7;
            14'd14850: out = 14'h11A7;
            14'd14851: out = 14'h11A7;
            14'd14852: out = 14'h11A7;
            14'd14853: out = 14'h11A6;
            14'd14854: out = 14'h11A6;
            14'd14855: out = 14'h11A6;
            14'd14856: out = 14'h11A5;
            14'd14857: out = 14'h11A5;
            14'd14858: out = 14'h11A5;
            14'd14859: out = 14'h11A4;
            14'd14860: out = 14'h11A4;
            14'd14861: out = 14'h11A4;
            14'd14862: out = 14'h11A3;
            14'd14863: out = 14'h11A3;
            14'd14864: out = 14'h11A3;
            14'd14865: out = 14'h11A3;
            14'd14866: out = 14'h11A2;
            14'd14867: out = 14'h11A2;
            14'd14868: out = 14'h11A2;
            14'd14869: out = 14'h11A1;
            14'd14870: out = 14'h11A1;
            14'd14871: out = 14'h11A1;
            14'd14872: out = 14'h11A0;
            14'd14873: out = 14'h11A0;
            14'd14874: out = 14'h11A0;
            14'd14875: out = 14'h11A0;
            14'd14876: out = 14'h119F;
            14'd14877: out = 14'h119F;
            14'd14878: out = 14'h119F;
            14'd14879: out = 14'h119E;
            14'd14880: out = 14'h119E;
            14'd14881: out = 14'h119E;
            14'd14882: out = 14'h119D;
            14'd14883: out = 14'h119D;
            14'd14884: out = 14'h119D;
            14'd14885: out = 14'h119C;
            14'd14886: out = 14'h119C;
            14'd14887: out = 14'h119C;
            14'd14888: out = 14'h119C;
            14'd14889: out = 14'h119B;
            14'd14890: out = 14'h119B;
            14'd14891: out = 14'h119B;
            14'd14892: out = 14'h119A;
            14'd14893: out = 14'h119A;
            14'd14894: out = 14'h119A;
            14'd14895: out = 14'h1199;
            14'd14896: out = 14'h1199;
            14'd14897: out = 14'h1199;
            14'd14898: out = 14'h1199;
            14'd14899: out = 14'h1198;
            14'd14900: out = 14'h1198;
            14'd14901: out = 14'h1198;
            14'd14902: out = 14'h1197;
            14'd14903: out = 14'h1197;
            14'd14904: out = 14'h1197;
            14'd14905: out = 14'h1196;
            14'd14906: out = 14'h1196;
            14'd14907: out = 14'h1196;
            14'd14908: out = 14'h1196;
            14'd14909: out = 14'h1195;
            14'd14910: out = 14'h1195;
            14'd14911: out = 14'h1195;
            14'd14912: out = 14'h1194;
            14'd14913: out = 14'h1194;
            14'd14914: out = 14'h1194;
            14'd14915: out = 14'h1193;
            14'd14916: out = 14'h1193;
            14'd14917: out = 14'h1193;
            14'd14918: out = 14'h1193;
            14'd14919: out = 14'h1192;
            14'd14920: out = 14'h1192;
            14'd14921: out = 14'h1192;
            14'd14922: out = 14'h1191;
            14'd14923: out = 14'h1191;
            14'd14924: out = 14'h1191;
            14'd14925: out = 14'h1190;
            14'd14926: out = 14'h1190;
            14'd14927: out = 14'h1190;
            14'd14928: out = 14'h1190;
            14'd14929: out = 14'h118F;
            14'd14930: out = 14'h118F;
            14'd14931: out = 14'h118F;
            14'd14932: out = 14'h118E;
            14'd14933: out = 14'h118E;
            14'd14934: out = 14'h118E;
            14'd14935: out = 14'h118D;
            14'd14936: out = 14'h118D;
            14'd14937: out = 14'h118D;
            14'd14938: out = 14'h118C;
            14'd14939: out = 14'h118C;
            14'd14940: out = 14'h118C;
            14'd14941: out = 14'h118C;
            14'd14942: out = 14'h118B;
            14'd14943: out = 14'h118B;
            14'd14944: out = 14'h118B;
            14'd14945: out = 14'h118A;
            14'd14946: out = 14'h118A;
            14'd14947: out = 14'h118A;
            14'd14948: out = 14'h1189;
            14'd14949: out = 14'h1189;
            14'd14950: out = 14'h1189;
            14'd14951: out = 14'h1189;
            14'd14952: out = 14'h1188;
            14'd14953: out = 14'h1188;
            14'd14954: out = 14'h1188;
            14'd14955: out = 14'h1187;
            14'd14956: out = 14'h1187;
            14'd14957: out = 14'h1187;
            14'd14958: out = 14'h1186;
            14'd14959: out = 14'h1186;
            14'd14960: out = 14'h1186;
            14'd14961: out = 14'h1186;
            14'd14962: out = 14'h1185;
            14'd14963: out = 14'h1185;
            14'd14964: out = 14'h1185;
            14'd14965: out = 14'h1184;
            14'd14966: out = 14'h1184;
            14'd14967: out = 14'h1184;
            14'd14968: out = 14'h1183;
            14'd14969: out = 14'h1183;
            14'd14970: out = 14'h1183;
            14'd14971: out = 14'h1183;
            14'd14972: out = 14'h1182;
            14'd14973: out = 14'h1182;
            14'd14974: out = 14'h1182;
            14'd14975: out = 14'h1181;
            14'd14976: out = 14'h1181;
            14'd14977: out = 14'h1181;
            14'd14978: out = 14'h1180;
            14'd14979: out = 14'h1180;
            14'd14980: out = 14'h1180;
            14'd14981: out = 14'h1180;
            14'd14982: out = 14'h117F;
            14'd14983: out = 14'h117F;
            14'd14984: out = 14'h117F;
            14'd14985: out = 14'h117E;
            14'd14986: out = 14'h117E;
            14'd14987: out = 14'h117E;
            14'd14988: out = 14'h117E;
            14'd14989: out = 14'h117D;
            14'd14990: out = 14'h117D;
            14'd14991: out = 14'h117D;
            14'd14992: out = 14'h117C;
            14'd14993: out = 14'h117C;
            14'd14994: out = 14'h117C;
            14'd14995: out = 14'h117B;
            14'd14996: out = 14'h117B;
            14'd14997: out = 14'h117B;
            14'd14998: out = 14'h117B;
            14'd14999: out = 14'h117A;
            14'd15000: out = 14'h117A;
            14'd15001: out = 14'h117A;
            14'd15002: out = 14'h1179;
            14'd15003: out = 14'h1179;
            14'd15004: out = 14'h1179;
            14'd15005: out = 14'h1178;
            14'd15006: out = 14'h1178;
            14'd15007: out = 14'h1178;
            14'd15008: out = 14'h1178;
            14'd15009: out = 14'h1177;
            14'd15010: out = 14'h1177;
            14'd15011: out = 14'h1177;
            14'd15012: out = 14'h1176;
            14'd15013: out = 14'h1176;
            14'd15014: out = 14'h1176;
            14'd15015: out = 14'h1175;
            14'd15016: out = 14'h1175;
            14'd15017: out = 14'h1175;
            14'd15018: out = 14'h1175;
            14'd15019: out = 14'h1174;
            14'd15020: out = 14'h1174;
            14'd15021: out = 14'h1174;
            14'd15022: out = 14'h1173;
            14'd15023: out = 14'h1173;
            14'd15024: out = 14'h1173;
            14'd15025: out = 14'h1172;
            14'd15026: out = 14'h1172;
            14'd15027: out = 14'h1172;
            14'd15028: out = 14'h1172;
            14'd15029: out = 14'h1171;
            14'd15030: out = 14'h1171;
            14'd15031: out = 14'h1171;
            14'd15032: out = 14'h1170;
            14'd15033: out = 14'h1170;
            14'd15034: out = 14'h1170;
            14'd15035: out = 14'h1170;
            14'd15036: out = 14'h116F;
            14'd15037: out = 14'h116F;
            14'd15038: out = 14'h116F;
            14'd15039: out = 14'h116E;
            14'd15040: out = 14'h116E;
            14'd15041: out = 14'h116E;
            14'd15042: out = 14'h116D;
            14'd15043: out = 14'h116D;
            14'd15044: out = 14'h116D;
            14'd15045: out = 14'h116D;
            14'd15046: out = 14'h116C;
            14'd15047: out = 14'h116C;
            14'd15048: out = 14'h116C;
            14'd15049: out = 14'h116B;
            14'd15050: out = 14'h116B;
            14'd15051: out = 14'h116B;
            14'd15052: out = 14'h116A;
            14'd15053: out = 14'h116A;
            14'd15054: out = 14'h116A;
            14'd15055: out = 14'h116A;
            14'd15056: out = 14'h1169;
            14'd15057: out = 14'h1169;
            14'd15058: out = 14'h1169;
            14'd15059: out = 14'h1168;
            14'd15060: out = 14'h1168;
            14'd15061: out = 14'h1168;
            14'd15062: out = 14'h1168;
            14'd15063: out = 14'h1167;
            14'd15064: out = 14'h1167;
            14'd15065: out = 14'h1167;
            14'd15066: out = 14'h1166;
            14'd15067: out = 14'h1166;
            14'd15068: out = 14'h1166;
            14'd15069: out = 14'h1165;
            14'd15070: out = 14'h1165;
            14'd15071: out = 14'h1165;
            14'd15072: out = 14'h1165;
            14'd15073: out = 14'h1164;
            14'd15074: out = 14'h1164;
            14'd15075: out = 14'h1164;
            14'd15076: out = 14'h1163;
            14'd15077: out = 14'h1163;
            14'd15078: out = 14'h1163;
            14'd15079: out = 14'h1162;
            14'd15080: out = 14'h1162;
            14'd15081: out = 14'h1162;
            14'd15082: out = 14'h1162;
            14'd15083: out = 14'h1161;
            14'd15084: out = 14'h1161;
            14'd15085: out = 14'h1161;
            14'd15086: out = 14'h1160;
            14'd15087: out = 14'h1160;
            14'd15088: out = 14'h1160;
            14'd15089: out = 14'h1160;
            14'd15090: out = 14'h115F;
            14'd15091: out = 14'h115F;
            14'd15092: out = 14'h115F;
            14'd15093: out = 14'h115E;
            14'd15094: out = 14'h115E;
            14'd15095: out = 14'h115E;
            14'd15096: out = 14'h115D;
            14'd15097: out = 14'h115D;
            14'd15098: out = 14'h115D;
            14'd15099: out = 14'h115D;
            14'd15100: out = 14'h115C;
            14'd15101: out = 14'h115C;
            14'd15102: out = 14'h115C;
            14'd15103: out = 14'h115B;
            14'd15104: out = 14'h115B;
            14'd15105: out = 14'h115B;
            14'd15106: out = 14'h115B;
            14'd15107: out = 14'h115A;
            14'd15108: out = 14'h115A;
            14'd15109: out = 14'h115A;
            14'd15110: out = 14'h1159;
            14'd15111: out = 14'h1159;
            14'd15112: out = 14'h1159;
            14'd15113: out = 14'h1158;
            14'd15114: out = 14'h1158;
            14'd15115: out = 14'h1158;
            14'd15116: out = 14'h1158;
            14'd15117: out = 14'h1157;
            14'd15118: out = 14'h1157;
            14'd15119: out = 14'h1157;
            14'd15120: out = 14'h1156;
            14'd15121: out = 14'h1156;
            14'd15122: out = 14'h1156;
            14'd15123: out = 14'h1156;
            14'd15124: out = 14'h1155;
            14'd15125: out = 14'h1155;
            14'd15126: out = 14'h1155;
            14'd15127: out = 14'h1154;
            14'd15128: out = 14'h1154;
            14'd15129: out = 14'h1154;
            14'd15130: out = 14'h1153;
            14'd15131: out = 14'h1153;
            14'd15132: out = 14'h1153;
            14'd15133: out = 14'h1153;
            14'd15134: out = 14'h1152;
            14'd15135: out = 14'h1152;
            14'd15136: out = 14'h1152;
            14'd15137: out = 14'h1151;
            14'd15138: out = 14'h1151;
            14'd15139: out = 14'h1151;
            14'd15140: out = 14'h1151;
            14'd15141: out = 14'h1150;
            14'd15142: out = 14'h1150;
            14'd15143: out = 14'h1150;
            14'd15144: out = 14'h114F;
            14'd15145: out = 14'h114F;
            14'd15146: out = 14'h114F;
            14'd15147: out = 14'h114F;
            14'd15148: out = 14'h114E;
            14'd15149: out = 14'h114E;
            14'd15150: out = 14'h114E;
            14'd15151: out = 14'h114D;
            14'd15152: out = 14'h114D;
            14'd15153: out = 14'h114D;
            14'd15154: out = 14'h114C;
            14'd15155: out = 14'h114C;
            14'd15156: out = 14'h114C;
            14'd15157: out = 14'h114C;
            14'd15158: out = 14'h114B;
            14'd15159: out = 14'h114B;
            14'd15160: out = 14'h114B;
            14'd15161: out = 14'h114A;
            14'd15162: out = 14'h114A;
            14'd15163: out = 14'h114A;
            14'd15164: out = 14'h114A;
            14'd15165: out = 14'h1149;
            14'd15166: out = 14'h1149;
            14'd15167: out = 14'h1149;
            14'd15168: out = 14'h1148;
            14'd15169: out = 14'h1148;
            14'd15170: out = 14'h1148;
            14'd15171: out = 14'h1147;
            14'd15172: out = 14'h1147;
            14'd15173: out = 14'h1147;
            14'd15174: out = 14'h1147;
            14'd15175: out = 14'h1146;
            14'd15176: out = 14'h1146;
            14'd15177: out = 14'h1146;
            14'd15178: out = 14'h1145;
            14'd15179: out = 14'h1145;
            14'd15180: out = 14'h1145;
            14'd15181: out = 14'h1145;
            14'd15182: out = 14'h1144;
            14'd15183: out = 14'h1144;
            14'd15184: out = 14'h1144;
            14'd15185: out = 14'h1143;
            14'd15186: out = 14'h1143;
            14'd15187: out = 14'h1143;
            14'd15188: out = 14'h1143;
            14'd15189: out = 14'h1142;
            14'd15190: out = 14'h1142;
            14'd15191: out = 14'h1142;
            14'd15192: out = 14'h1141;
            14'd15193: out = 14'h1141;
            14'd15194: out = 14'h1141;
            14'd15195: out = 14'h1141;
            14'd15196: out = 14'h1140;
            14'd15197: out = 14'h1140;
            14'd15198: out = 14'h1140;
            14'd15199: out = 14'h113F;
            14'd15200: out = 14'h113F;
            14'd15201: out = 14'h113F;
            14'd15202: out = 14'h113E;
            14'd15203: out = 14'h113E;
            14'd15204: out = 14'h113E;
            14'd15205: out = 14'h113E;
            14'd15206: out = 14'h113D;
            14'd15207: out = 14'h113D;
            14'd15208: out = 14'h113D;
            14'd15209: out = 14'h113C;
            14'd15210: out = 14'h113C;
            14'd15211: out = 14'h113C;
            14'd15212: out = 14'h113C;
            14'd15213: out = 14'h113B;
            14'd15214: out = 14'h113B;
            14'd15215: out = 14'h113B;
            14'd15216: out = 14'h113A;
            14'd15217: out = 14'h113A;
            14'd15218: out = 14'h113A;
            14'd15219: out = 14'h113A;
            14'd15220: out = 14'h1139;
            14'd15221: out = 14'h1139;
            14'd15222: out = 14'h1139;
            14'd15223: out = 14'h1138;
            14'd15224: out = 14'h1138;
            14'd15225: out = 14'h1138;
            14'd15226: out = 14'h1138;
            14'd15227: out = 14'h1137;
            14'd15228: out = 14'h1137;
            14'd15229: out = 14'h1137;
            14'd15230: out = 14'h1136;
            14'd15231: out = 14'h1136;
            14'd15232: out = 14'h1136;
            14'd15233: out = 14'h1135;
            14'd15234: out = 14'h1135;
            14'd15235: out = 14'h1135;
            14'd15236: out = 14'h1135;
            14'd15237: out = 14'h1134;
            14'd15238: out = 14'h1134;
            14'd15239: out = 14'h1134;
            14'd15240: out = 14'h1133;
            14'd15241: out = 14'h1133;
            14'd15242: out = 14'h1133;
            14'd15243: out = 14'h1133;
            14'd15244: out = 14'h1132;
            14'd15245: out = 14'h1132;
            14'd15246: out = 14'h1132;
            14'd15247: out = 14'h1131;
            14'd15248: out = 14'h1131;
            14'd15249: out = 14'h1131;
            14'd15250: out = 14'h1131;
            14'd15251: out = 14'h1130;
            14'd15252: out = 14'h1130;
            14'd15253: out = 14'h1130;
            14'd15254: out = 14'h112F;
            14'd15255: out = 14'h112F;
            14'd15256: out = 14'h112F;
            14'd15257: out = 14'h112F;
            14'd15258: out = 14'h112E;
            14'd15259: out = 14'h112E;
            14'd15260: out = 14'h112E;
            14'd15261: out = 14'h112D;
            14'd15262: out = 14'h112D;
            14'd15263: out = 14'h112D;
            14'd15264: out = 14'h112D;
            14'd15265: out = 14'h112C;
            14'd15266: out = 14'h112C;
            14'd15267: out = 14'h112C;
            14'd15268: out = 14'h112B;
            14'd15269: out = 14'h112B;
            14'd15270: out = 14'h112B;
            14'd15271: out = 14'h112B;
            14'd15272: out = 14'h112A;
            14'd15273: out = 14'h112A;
            14'd15274: out = 14'h112A;
            14'd15275: out = 14'h1129;
            14'd15276: out = 14'h1129;
            14'd15277: out = 14'h1129;
            14'd15278: out = 14'h1129;
            14'd15279: out = 14'h1128;
            14'd15280: out = 14'h1128;
            14'd15281: out = 14'h1128;
            14'd15282: out = 14'h1127;
            14'd15283: out = 14'h1127;
            14'd15284: out = 14'h1127;
            14'd15285: out = 14'h1127;
            14'd15286: out = 14'h1126;
            14'd15287: out = 14'h1126;
            14'd15288: out = 14'h1126;
            14'd15289: out = 14'h1125;
            14'd15290: out = 14'h1125;
            14'd15291: out = 14'h1125;
            14'd15292: out = 14'h1124;
            14'd15293: out = 14'h1124;
            14'd15294: out = 14'h1124;
            14'd15295: out = 14'h1124;
            14'd15296: out = 14'h1123;
            14'd15297: out = 14'h1123;
            14'd15298: out = 14'h1123;
            14'd15299: out = 14'h1122;
            14'd15300: out = 14'h1122;
            14'd15301: out = 14'h1122;
            14'd15302: out = 14'h1122;
            14'd15303: out = 14'h1121;
            14'd15304: out = 14'h1121;
            14'd15305: out = 14'h1121;
            14'd15306: out = 14'h1120;
            14'd15307: out = 14'h1120;
            14'd15308: out = 14'h1120;
            14'd15309: out = 14'h1120;
            14'd15310: out = 14'h111F;
            14'd15311: out = 14'h111F;
            14'd15312: out = 14'h111F;
            14'd15313: out = 14'h111E;
            14'd15314: out = 14'h111E;
            14'd15315: out = 14'h111E;
            14'd15316: out = 14'h111E;
            14'd15317: out = 14'h111D;
            14'd15318: out = 14'h111D;
            14'd15319: out = 14'h111D;
            14'd15320: out = 14'h111C;
            14'd15321: out = 14'h111C;
            14'd15322: out = 14'h111C;
            14'd15323: out = 14'h111C;
            14'd15324: out = 14'h111B;
            14'd15325: out = 14'h111B;
            14'd15326: out = 14'h111B;
            14'd15327: out = 14'h111A;
            14'd15328: out = 14'h111A;
            14'd15329: out = 14'h111A;
            14'd15330: out = 14'h111A;
            14'd15331: out = 14'h1119;
            14'd15332: out = 14'h1119;
            14'd15333: out = 14'h1119;
            14'd15334: out = 14'h1118;
            14'd15335: out = 14'h1118;
            14'd15336: out = 14'h1118;
            14'd15337: out = 14'h1118;
            14'd15338: out = 14'h1117;
            14'd15339: out = 14'h1117;
            14'd15340: out = 14'h1117;
            14'd15341: out = 14'h1116;
            14'd15342: out = 14'h1116;
            14'd15343: out = 14'h1116;
            14'd15344: out = 14'h1116;
            14'd15345: out = 14'h1115;
            14'd15346: out = 14'h1115;
            14'd15347: out = 14'h1115;
            14'd15348: out = 14'h1114;
            14'd15349: out = 14'h1114;
            14'd15350: out = 14'h1114;
            14'd15351: out = 14'h1114;
            14'd15352: out = 14'h1113;
            14'd15353: out = 14'h1113;
            14'd15354: out = 14'h1113;
            14'd15355: out = 14'h1112;
            14'd15356: out = 14'h1112;
            14'd15357: out = 14'h1112;
            14'd15358: out = 14'h1112;
            14'd15359: out = 14'h1111;
            14'd15360: out = 14'h1111;
            14'd15361: out = 14'h1111;
            14'd15362: out = 14'h1110;
            14'd15363: out = 14'h1110;
            14'd15364: out = 14'h1110;
            14'd15365: out = 14'h1110;
            14'd15366: out = 14'h110F;
            14'd15367: out = 14'h110F;
            14'd15368: out = 14'h110F;
            14'd15369: out = 14'h110F;
            14'd15370: out = 14'h110E;
            14'd15371: out = 14'h110E;
            14'd15372: out = 14'h110E;
            14'd15373: out = 14'h110D;
            14'd15374: out = 14'h110D;
            14'd15375: out = 14'h110D;
            14'd15376: out = 14'h110D;
            14'd15377: out = 14'h110C;
            14'd15378: out = 14'h110C;
            14'd15379: out = 14'h110C;
            14'd15380: out = 14'h110B;
            14'd15381: out = 14'h110B;
            14'd15382: out = 14'h110B;
            14'd15383: out = 14'h110B;
            14'd15384: out = 14'h110A;
            14'd15385: out = 14'h110A;
            14'd15386: out = 14'h110A;
            14'd15387: out = 14'h1109;
            14'd15388: out = 14'h1109;
            14'd15389: out = 14'h1109;
            14'd15390: out = 14'h1109;
            14'd15391: out = 14'h1108;
            14'd15392: out = 14'h1108;
            14'd15393: out = 14'h1108;
            14'd15394: out = 14'h1107;
            14'd15395: out = 14'h1107;
            14'd15396: out = 14'h1107;
            14'd15397: out = 14'h1107;
            14'd15398: out = 14'h1106;
            14'd15399: out = 14'h1106;
            14'd15400: out = 14'h1106;
            14'd15401: out = 14'h1105;
            14'd15402: out = 14'h1105;
            14'd15403: out = 14'h1105;
            14'd15404: out = 14'h1105;
            14'd15405: out = 14'h1104;
            14'd15406: out = 14'h1104;
            14'd15407: out = 14'h1104;
            14'd15408: out = 14'h1103;
            14'd15409: out = 14'h1103;
            14'd15410: out = 14'h1103;
            14'd15411: out = 14'h1103;
            14'd15412: out = 14'h1102;
            14'd15413: out = 14'h1102;
            14'd15414: out = 14'h1102;
            14'd15415: out = 14'h1101;
            14'd15416: out = 14'h1101;
            14'd15417: out = 14'h1101;
            14'd15418: out = 14'h1101;
            14'd15419: out = 14'h1100;
            14'd15420: out = 14'h1100;
            14'd15421: out = 14'h1100;
            14'd15422: out = 14'h1100;
            14'd15423: out = 14'h10FF;
            14'd15424: out = 14'h10FF;
            14'd15425: out = 14'h10FF;
            14'd15426: out = 14'h10FE;
            14'd15427: out = 14'h10FE;
            14'd15428: out = 14'h10FE;
            14'd15429: out = 14'h10FE;
            14'd15430: out = 14'h10FD;
            14'd15431: out = 14'h10FD;
            14'd15432: out = 14'h10FD;
            14'd15433: out = 14'h10FC;
            14'd15434: out = 14'h10FC;
            14'd15435: out = 14'h10FC;
            14'd15436: out = 14'h10FC;
            14'd15437: out = 14'h10FB;
            14'd15438: out = 14'h10FB;
            14'd15439: out = 14'h10FB;
            14'd15440: out = 14'h10FA;
            14'd15441: out = 14'h10FA;
            14'd15442: out = 14'h10FA;
            14'd15443: out = 14'h10FA;
            14'd15444: out = 14'h10F9;
            14'd15445: out = 14'h10F9;
            14'd15446: out = 14'h10F9;
            14'd15447: out = 14'h10F8;
            14'd15448: out = 14'h10F8;
            14'd15449: out = 14'h10F8;
            14'd15450: out = 14'h10F8;
            14'd15451: out = 14'h10F7;
            14'd15452: out = 14'h10F7;
            14'd15453: out = 14'h10F7;
            14'd15454: out = 14'h10F6;
            14'd15455: out = 14'h10F6;
            14'd15456: out = 14'h10F6;
            14'd15457: out = 14'h10F6;
            14'd15458: out = 14'h10F5;
            14'd15459: out = 14'h10F5;
            14'd15460: out = 14'h10F5;
            14'd15461: out = 14'h10F5;
            14'd15462: out = 14'h10F4;
            14'd15463: out = 14'h10F4;
            14'd15464: out = 14'h10F4;
            14'd15465: out = 14'h10F3;
            14'd15466: out = 14'h10F3;
            14'd15467: out = 14'h10F3;
            14'd15468: out = 14'h10F3;
            14'd15469: out = 14'h10F2;
            14'd15470: out = 14'h10F2;
            14'd15471: out = 14'h10F2;
            14'd15472: out = 14'h10F1;
            14'd15473: out = 14'h10F1;
            14'd15474: out = 14'h10F1;
            14'd15475: out = 14'h10F1;
            14'd15476: out = 14'h10F0;
            14'd15477: out = 14'h10F0;
            14'd15478: out = 14'h10F0;
            14'd15479: out = 14'h10EF;
            14'd15480: out = 14'h10EF;
            14'd15481: out = 14'h10EF;
            14'd15482: out = 14'h10EF;
            14'd15483: out = 14'h10EE;
            14'd15484: out = 14'h10EE;
            14'd15485: out = 14'h10EE;
            14'd15486: out = 14'h10EE;
            14'd15487: out = 14'h10ED;
            14'd15488: out = 14'h10ED;
            14'd15489: out = 14'h10ED;
            14'd15490: out = 14'h10EC;
            14'd15491: out = 14'h10EC;
            14'd15492: out = 14'h10EC;
            14'd15493: out = 14'h10EC;
            14'd15494: out = 14'h10EB;
            14'd15495: out = 14'h10EB;
            14'd15496: out = 14'h10EB;
            14'd15497: out = 14'h10EA;
            14'd15498: out = 14'h10EA;
            14'd15499: out = 14'h10EA;
            14'd15500: out = 14'h10EA;
            14'd15501: out = 14'h10E9;
            14'd15502: out = 14'h10E9;
            14'd15503: out = 14'h10E9;
            14'd15504: out = 14'h10E8;
            14'd15505: out = 14'h10E8;
            14'd15506: out = 14'h10E8;
            14'd15507: out = 14'h10E8;
            14'd15508: out = 14'h10E7;
            14'd15509: out = 14'h10E7;
            14'd15510: out = 14'h10E7;
            14'd15511: out = 14'h10E7;
            14'd15512: out = 14'h10E6;
            14'd15513: out = 14'h10E6;
            14'd15514: out = 14'h10E6;
            14'd15515: out = 14'h10E5;
            14'd15516: out = 14'h10E5;
            14'd15517: out = 14'h10E5;
            14'd15518: out = 14'h10E5;
            14'd15519: out = 14'h10E4;
            14'd15520: out = 14'h10E4;
            14'd15521: out = 14'h10E4;
            14'd15522: out = 14'h10E3;
            14'd15523: out = 14'h10E3;
            14'd15524: out = 14'h10E3;
            14'd15525: out = 14'h10E3;
            14'd15526: out = 14'h10E2;
            14'd15527: out = 14'h10E2;
            14'd15528: out = 14'h10E2;
            14'd15529: out = 14'h10E2;
            14'd15530: out = 14'h10E1;
            14'd15531: out = 14'h10E1;
            14'd15532: out = 14'h10E1;
            14'd15533: out = 14'h10E0;
            14'd15534: out = 14'h10E0;
            14'd15535: out = 14'h10E0;
            14'd15536: out = 14'h10E0;
            14'd15537: out = 14'h10DF;
            14'd15538: out = 14'h10DF;
            14'd15539: out = 14'h10DF;
            14'd15540: out = 14'h10DE;
            14'd15541: out = 14'h10DE;
            14'd15542: out = 14'h10DE;
            14'd15543: out = 14'h10DE;
            14'd15544: out = 14'h10DD;
            14'd15545: out = 14'h10DD;
            14'd15546: out = 14'h10DD;
            14'd15547: out = 14'h10DD;
            14'd15548: out = 14'h10DC;
            14'd15549: out = 14'h10DC;
            14'd15550: out = 14'h10DC;
            14'd15551: out = 14'h10DB;
            14'd15552: out = 14'h10DB;
            14'd15553: out = 14'h10DB;
            14'd15554: out = 14'h10DB;
            14'd15555: out = 14'h10DA;
            14'd15556: out = 14'h10DA;
            14'd15557: out = 14'h10DA;
            14'd15558: out = 14'h10D9;
            14'd15559: out = 14'h10D9;
            14'd15560: out = 14'h10D9;
            14'd15561: out = 14'h10D9;
            14'd15562: out = 14'h10D8;
            14'd15563: out = 14'h10D8;
            14'd15564: out = 14'h10D8;
            14'd15565: out = 14'h10D8;
            14'd15566: out = 14'h10D7;
            14'd15567: out = 14'h10D7;
            14'd15568: out = 14'h10D7;
            14'd15569: out = 14'h10D6;
            14'd15570: out = 14'h10D6;
            14'd15571: out = 14'h10D6;
            14'd15572: out = 14'h10D6;
            14'd15573: out = 14'h10D5;
            14'd15574: out = 14'h10D5;
            14'd15575: out = 14'h10D5;
            14'd15576: out = 14'h10D4;
            14'd15577: out = 14'h10D4;
            14'd15578: out = 14'h10D4;
            14'd15579: out = 14'h10D4;
            14'd15580: out = 14'h10D3;
            14'd15581: out = 14'h10D3;
            14'd15582: out = 14'h10D3;
            14'd15583: out = 14'h10D3;
            14'd15584: out = 14'h10D2;
            14'd15585: out = 14'h10D2;
            14'd15586: out = 14'h10D2;
            14'd15587: out = 14'h10D1;
            14'd15588: out = 14'h10D1;
            14'd15589: out = 14'h10D1;
            14'd15590: out = 14'h10D1;
            14'd15591: out = 14'h10D0;
            14'd15592: out = 14'h10D0;
            14'd15593: out = 14'h10D0;
            14'd15594: out = 14'h10D0;
            14'd15595: out = 14'h10CF;
            14'd15596: out = 14'h10CF;
            14'd15597: out = 14'h10CF;
            14'd15598: out = 14'h10CE;
            14'd15599: out = 14'h10CE;
            14'd15600: out = 14'h10CE;
            14'd15601: out = 14'h10CE;
            14'd15602: out = 14'h10CD;
            14'd15603: out = 14'h10CD;
            14'd15604: out = 14'h10CD;
            14'd15605: out = 14'h10CC;
            14'd15606: out = 14'h10CC;
            14'd15607: out = 14'h10CC;
            14'd15608: out = 14'h10CC;
            14'd15609: out = 14'h10CB;
            14'd15610: out = 14'h10CB;
            14'd15611: out = 14'h10CB;
            14'd15612: out = 14'h10CB;
            14'd15613: out = 14'h10CA;
            14'd15614: out = 14'h10CA;
            14'd15615: out = 14'h10CA;
            14'd15616: out = 14'h10C9;
            14'd15617: out = 14'h10C9;
            14'd15618: out = 14'h10C9;
            14'd15619: out = 14'h10C9;
            14'd15620: out = 14'h10C8;
            14'd15621: out = 14'h10C8;
            14'd15622: out = 14'h10C8;
            14'd15623: out = 14'h10C8;
            14'd15624: out = 14'h10C7;
            14'd15625: out = 14'h10C7;
            14'd15626: out = 14'h10C7;
            14'd15627: out = 14'h10C6;
            14'd15628: out = 14'h10C6;
            14'd15629: out = 14'h10C6;
            14'd15630: out = 14'h10C6;
            14'd15631: out = 14'h10C5;
            14'd15632: out = 14'h10C5;
            14'd15633: out = 14'h10C5;
            14'd15634: out = 14'h10C4;
            14'd15635: out = 14'h10C4;
            14'd15636: out = 14'h10C4;
            14'd15637: out = 14'h10C4;
            14'd15638: out = 14'h10C3;
            14'd15639: out = 14'h10C3;
            14'd15640: out = 14'h10C3;
            14'd15641: out = 14'h10C3;
            14'd15642: out = 14'h10C2;
            14'd15643: out = 14'h10C2;
            14'd15644: out = 14'h10C2;
            14'd15645: out = 14'h10C1;
            14'd15646: out = 14'h10C1;
            14'd15647: out = 14'h10C1;
            14'd15648: out = 14'h10C1;
            14'd15649: out = 14'h10C0;
            14'd15650: out = 14'h10C0;
            14'd15651: out = 14'h10C0;
            14'd15652: out = 14'h10C0;
            14'd15653: out = 14'h10BF;
            14'd15654: out = 14'h10BF;
            14'd15655: out = 14'h10BF;
            14'd15656: out = 14'h10BE;
            14'd15657: out = 14'h10BE;
            14'd15658: out = 14'h10BE;
            14'd15659: out = 14'h10BE;
            14'd15660: out = 14'h10BD;
            14'd15661: out = 14'h10BD;
            14'd15662: out = 14'h10BD;
            14'd15663: out = 14'h10BD;
            14'd15664: out = 14'h10BC;
            14'd15665: out = 14'h10BC;
            14'd15666: out = 14'h10BC;
            14'd15667: out = 14'h10BB;
            14'd15668: out = 14'h10BB;
            14'd15669: out = 14'h10BB;
            14'd15670: out = 14'h10BB;
            14'd15671: out = 14'h10BA;
            14'd15672: out = 14'h10BA;
            14'd15673: out = 14'h10BA;
            14'd15674: out = 14'h10BA;
            14'd15675: out = 14'h10B9;
            14'd15676: out = 14'h10B9;
            14'd15677: out = 14'h10B9;
            14'd15678: out = 14'h10B8;
            14'd15679: out = 14'h10B8;
            14'd15680: out = 14'h10B8;
            14'd15681: out = 14'h10B8;
            14'd15682: out = 14'h10B7;
            14'd15683: out = 14'h10B7;
            14'd15684: out = 14'h10B7;
            14'd15685: out = 14'h10B7;
            14'd15686: out = 14'h10B6;
            14'd15687: out = 14'h10B6;
            14'd15688: out = 14'h10B6;
            14'd15689: out = 14'h10B5;
            14'd15690: out = 14'h10B5;
            14'd15691: out = 14'h10B5;
            14'd15692: out = 14'h10B5;
            14'd15693: out = 14'h10B4;
            14'd15694: out = 14'h10B4;
            14'd15695: out = 14'h10B4;
            14'd15696: out = 14'h10B4;
            14'd15697: out = 14'h10B3;
            14'd15698: out = 14'h10B3;
            14'd15699: out = 14'h10B3;
            14'd15700: out = 14'h10B2;
            14'd15701: out = 14'h10B2;
            14'd15702: out = 14'h10B2;
            14'd15703: out = 14'h10B2;
            14'd15704: out = 14'h10B1;
            14'd15705: out = 14'h10B1;
            14'd15706: out = 14'h10B1;
            14'd15707: out = 14'h10B1;
            14'd15708: out = 14'h10B0;
            14'd15709: out = 14'h10B0;
            14'd15710: out = 14'h10B0;
            14'd15711: out = 14'h10AF;
            14'd15712: out = 14'h10AF;
            14'd15713: out = 14'h10AF;
            14'd15714: out = 14'h10AF;
            14'd15715: out = 14'h10AE;
            14'd15716: out = 14'h10AE;
            14'd15717: out = 14'h10AE;
            14'd15718: out = 14'h10AE;
            14'd15719: out = 14'h10AD;
            14'd15720: out = 14'h10AD;
            14'd15721: out = 14'h10AD;
            14'd15722: out = 14'h10AC;
            14'd15723: out = 14'h10AC;
            14'd15724: out = 14'h10AC;
            14'd15725: out = 14'h10AC;
            14'd15726: out = 14'h10AB;
            14'd15727: out = 14'h10AB;
            14'd15728: out = 14'h10AB;
            14'd15729: out = 14'h10AB;
            14'd15730: out = 14'h10AA;
            14'd15731: out = 14'h10AA;
            14'd15732: out = 14'h10AA;
            14'd15733: out = 14'h10A9;
            14'd15734: out = 14'h10A9;
            14'd15735: out = 14'h10A9;
            14'd15736: out = 14'h10A9;
            14'd15737: out = 14'h10A8;
            14'd15738: out = 14'h10A8;
            14'd15739: out = 14'h10A8;
            14'd15740: out = 14'h10A8;
            14'd15741: out = 14'h10A7;
            14'd15742: out = 14'h10A7;
            14'd15743: out = 14'h10A7;
            14'd15744: out = 14'h10A7;
            14'd15745: out = 14'h10A6;
            14'd15746: out = 14'h10A6;
            14'd15747: out = 14'h10A6;
            14'd15748: out = 14'h10A5;
            14'd15749: out = 14'h10A5;
            14'd15750: out = 14'h10A5;
            14'd15751: out = 14'h10A5;
            14'd15752: out = 14'h10A4;
            14'd15753: out = 14'h10A4;
            14'd15754: out = 14'h10A4;
            14'd15755: out = 14'h10A4;
            14'd15756: out = 14'h10A3;
            14'd15757: out = 14'h10A3;
            14'd15758: out = 14'h10A3;
            14'd15759: out = 14'h10A2;
            14'd15760: out = 14'h10A2;
            14'd15761: out = 14'h10A2;
            14'd15762: out = 14'h10A2;
            14'd15763: out = 14'h10A1;
            14'd15764: out = 14'h10A1;
            14'd15765: out = 14'h10A1;
            14'd15766: out = 14'h10A1;
            14'd15767: out = 14'h10A0;
            14'd15768: out = 14'h10A0;
            14'd15769: out = 14'h10A0;
            14'd15770: out = 14'h109F;
            14'd15771: out = 14'h109F;
            14'd15772: out = 14'h109F;
            14'd15773: out = 14'h109F;
            14'd15774: out = 14'h109E;
            14'd15775: out = 14'h109E;
            14'd15776: out = 14'h109E;
            14'd15777: out = 14'h109E;
            14'd15778: out = 14'h109D;
            14'd15779: out = 14'h109D;
            14'd15780: out = 14'h109D;
            14'd15781: out = 14'h109D;
            14'd15782: out = 14'h109C;
            14'd15783: out = 14'h109C;
            14'd15784: out = 14'h109C;
            14'd15785: out = 14'h109B;
            14'd15786: out = 14'h109B;
            14'd15787: out = 14'h109B;
            14'd15788: out = 14'h109B;
            14'd15789: out = 14'h109A;
            14'd15790: out = 14'h109A;
            14'd15791: out = 14'h109A;
            14'd15792: out = 14'h109A;
            14'd15793: out = 14'h1099;
            14'd15794: out = 14'h1099;
            14'd15795: out = 14'h1099;
            14'd15796: out = 14'h1098;
            14'd15797: out = 14'h1098;
            14'd15798: out = 14'h1098;
            14'd15799: out = 14'h1098;
            14'd15800: out = 14'h1097;
            14'd15801: out = 14'h1097;
            14'd15802: out = 14'h1097;
            14'd15803: out = 14'h1097;
            14'd15804: out = 14'h1096;
            14'd15805: out = 14'h1096;
            14'd15806: out = 14'h1096;
            14'd15807: out = 14'h1096;
            14'd15808: out = 14'h1095;
            14'd15809: out = 14'h1095;
            14'd15810: out = 14'h1095;
            14'd15811: out = 14'h1094;
            14'd15812: out = 14'h1094;
            14'd15813: out = 14'h1094;
            14'd15814: out = 14'h1094;
            14'd15815: out = 14'h1093;
            14'd15816: out = 14'h1093;
            14'd15817: out = 14'h1093;
            14'd15818: out = 14'h1093;
            14'd15819: out = 14'h1092;
            14'd15820: out = 14'h1092;
            14'd15821: out = 14'h1092;
            14'd15822: out = 14'h1091;
            14'd15823: out = 14'h1091;
            14'd15824: out = 14'h1091;
            14'd15825: out = 14'h1091;
            14'd15826: out = 14'h1090;
            14'd15827: out = 14'h1090;
            14'd15828: out = 14'h1090;
            14'd15829: out = 14'h1090;
            14'd15830: out = 14'h108F;
            14'd15831: out = 14'h108F;
            14'd15832: out = 14'h108F;
            14'd15833: out = 14'h108F;
            14'd15834: out = 14'h108E;
            14'd15835: out = 14'h108E;
            14'd15836: out = 14'h108E;
            14'd15837: out = 14'h108D;
            14'd15838: out = 14'h108D;
            14'd15839: out = 14'h108D;
            14'd15840: out = 14'h108D;
            14'd15841: out = 14'h108C;
            14'd15842: out = 14'h108C;
            14'd15843: out = 14'h108C;
            14'd15844: out = 14'h108C;
            14'd15845: out = 14'h108B;
            14'd15846: out = 14'h108B;
            14'd15847: out = 14'h108B;
            14'd15848: out = 14'h108B;
            14'd15849: out = 14'h108A;
            14'd15850: out = 14'h108A;
            14'd15851: out = 14'h108A;
            14'd15852: out = 14'h1089;
            14'd15853: out = 14'h1089;
            14'd15854: out = 14'h1089;
            14'd15855: out = 14'h1089;
            14'd15856: out = 14'h1088;
            14'd15857: out = 14'h1088;
            14'd15858: out = 14'h1088;
            14'd15859: out = 14'h1088;
            14'd15860: out = 14'h1087;
            14'd15861: out = 14'h1087;
            14'd15862: out = 14'h1087;
            14'd15863: out = 14'h1087;
            14'd15864: out = 14'h1086;
            14'd15865: out = 14'h1086;
            14'd15866: out = 14'h1086;
            14'd15867: out = 14'h1085;
            14'd15868: out = 14'h1085;
            14'd15869: out = 14'h1085;
            14'd15870: out = 14'h1085;
            14'd15871: out = 14'h1084;
            14'd15872: out = 14'h1084;
            14'd15873: out = 14'h1084;
            14'd15874: out = 14'h1084;
            14'd15875: out = 14'h1083;
            14'd15876: out = 14'h1083;
            14'd15877: out = 14'h1083;
            14'd15878: out = 14'h1083;
            14'd15879: out = 14'h1082;
            14'd15880: out = 14'h1082;
            14'd15881: out = 14'h1082;
            14'd15882: out = 14'h1081;
            14'd15883: out = 14'h1081;
            14'd15884: out = 14'h1081;
            14'd15885: out = 14'h1081;
            14'd15886: out = 14'h1080;
            14'd15887: out = 14'h1080;
            14'd15888: out = 14'h1080;
            14'd15889: out = 14'h1080;
            14'd15890: out = 14'h107F;
            14'd15891: out = 14'h107F;
            14'd15892: out = 14'h107F;
            14'd15893: out = 14'h107F;
            14'd15894: out = 14'h107E;
            14'd15895: out = 14'h107E;
            14'd15896: out = 14'h107E;
            14'd15897: out = 14'h107D;
            14'd15898: out = 14'h107D;
            14'd15899: out = 14'h107D;
            14'd15900: out = 14'h107D;
            14'd15901: out = 14'h107C;
            14'd15902: out = 14'h107C;
            14'd15903: out = 14'h107C;
            14'd15904: out = 14'h107C;
            14'd15905: out = 14'h107B;
            14'd15906: out = 14'h107B;
            14'd15907: out = 14'h107B;
            14'd15908: out = 14'h107B;
            14'd15909: out = 14'h107A;
            14'd15910: out = 14'h107A;
            14'd15911: out = 14'h107A;
            14'd15912: out = 14'h107A;
            14'd15913: out = 14'h1079;
            14'd15914: out = 14'h1079;
            14'd15915: out = 14'h1079;
            14'd15916: out = 14'h1078;
            14'd15917: out = 14'h1078;
            14'd15918: out = 14'h1078;
            14'd15919: out = 14'h1078;
            14'd15920: out = 14'h1077;
            14'd15921: out = 14'h1077;
            14'd15922: out = 14'h1077;
            14'd15923: out = 14'h1077;
            14'd15924: out = 14'h1076;
            14'd15925: out = 14'h1076;
            14'd15926: out = 14'h1076;
            14'd15927: out = 14'h1076;
            14'd15928: out = 14'h1075;
            14'd15929: out = 14'h1075;
            14'd15930: out = 14'h1075;
            14'd15931: out = 14'h1074;
            14'd15932: out = 14'h1074;
            14'd15933: out = 14'h1074;
            14'd15934: out = 14'h1074;
            14'd15935: out = 14'h1073;
            14'd15936: out = 14'h1073;
            14'd15937: out = 14'h1073;
            14'd15938: out = 14'h1073;
            14'd15939: out = 14'h1072;
            14'd15940: out = 14'h1072;
            14'd15941: out = 14'h1072;
            14'd15942: out = 14'h1072;
            14'd15943: out = 14'h1071;
            14'd15944: out = 14'h1071;
            14'd15945: out = 14'h1071;
            14'd15946: out = 14'h1071;
            14'd15947: out = 14'h1070;
            14'd15948: out = 14'h1070;
            14'd15949: out = 14'h1070;
            14'd15950: out = 14'h106F;
            14'd15951: out = 14'h106F;
            14'd15952: out = 14'h106F;
            14'd15953: out = 14'h106F;
            14'd15954: out = 14'h106E;
            14'd15955: out = 14'h106E;
            14'd15956: out = 14'h106E;
            14'd15957: out = 14'h106E;
            14'd15958: out = 14'h106D;
            14'd15959: out = 14'h106D;
            14'd15960: out = 14'h106D;
            14'd15961: out = 14'h106D;
            14'd15962: out = 14'h106C;
            14'd15963: out = 14'h106C;
            14'd15964: out = 14'h106C;
            14'd15965: out = 14'h106B;
            14'd15966: out = 14'h106B;
            14'd15967: out = 14'h106B;
            14'd15968: out = 14'h106B;
            14'd15969: out = 14'h106A;
            14'd15970: out = 14'h106A;
            14'd15971: out = 14'h106A;
            14'd15972: out = 14'h106A;
            14'd15973: out = 14'h1069;
            14'd15974: out = 14'h1069;
            14'd15975: out = 14'h1069;
            14'd15976: out = 14'h1069;
            14'd15977: out = 14'h1068;
            14'd15978: out = 14'h1068;
            14'd15979: out = 14'h1068;
            14'd15980: out = 14'h1068;
            14'd15981: out = 14'h1067;
            14'd15982: out = 14'h1067;
            14'd15983: out = 14'h1067;
            14'd15984: out = 14'h1067;
            14'd15985: out = 14'h1066;
            14'd15986: out = 14'h1066;
            14'd15987: out = 14'h1066;
            14'd15988: out = 14'h1065;
            14'd15989: out = 14'h1065;
            14'd15990: out = 14'h1065;
            14'd15991: out = 14'h1065;
            14'd15992: out = 14'h1064;
            14'd15993: out = 14'h1064;
            14'd15994: out = 14'h1064;
            14'd15995: out = 14'h1064;
            14'd15996: out = 14'h1063;
            14'd15997: out = 14'h1063;
            14'd15998: out = 14'h1063;
            14'd15999: out = 14'h1063;
            14'd16000: out = 14'h1062;
            14'd16001: out = 14'h1062;
            14'd16002: out = 14'h1062;
            14'd16003: out = 14'h1062;
            14'd16004: out = 14'h1061;
            14'd16005: out = 14'h1061;
            14'd16006: out = 14'h1061;
            14'd16007: out = 14'h1060;
            14'd16008: out = 14'h1060;
            14'd16009: out = 14'h1060;
            14'd16010: out = 14'h1060;
            14'd16011: out = 14'h105F;
            14'd16012: out = 14'h105F;
            14'd16013: out = 14'h105F;
            14'd16014: out = 14'h105F;
            14'd16015: out = 14'h105E;
            14'd16016: out = 14'h105E;
            14'd16017: out = 14'h105E;
            14'd16018: out = 14'h105E;
            14'd16019: out = 14'h105D;
            14'd16020: out = 14'h105D;
            14'd16021: out = 14'h105D;
            14'd16022: out = 14'h105D;
            14'd16023: out = 14'h105C;
            14'd16024: out = 14'h105C;
            14'd16025: out = 14'h105C;
            14'd16026: out = 14'h105B;
            14'd16027: out = 14'h105B;
            14'd16028: out = 14'h105B;
            14'd16029: out = 14'h105B;
            14'd16030: out = 14'h105A;
            14'd16031: out = 14'h105A;
            14'd16032: out = 14'h105A;
            14'd16033: out = 14'h105A;
            14'd16034: out = 14'h1059;
            14'd16035: out = 14'h1059;
            14'd16036: out = 14'h1059;
            14'd16037: out = 14'h1059;
            14'd16038: out = 14'h1058;
            14'd16039: out = 14'h1058;
            14'd16040: out = 14'h1058;
            14'd16041: out = 14'h1058;
            14'd16042: out = 14'h1057;
            14'd16043: out = 14'h1057;
            14'd16044: out = 14'h1057;
            14'd16045: out = 14'h1057;
            14'd16046: out = 14'h1056;
            14'd16047: out = 14'h1056;
            14'd16048: out = 14'h1056;
            14'd16049: out = 14'h1055;
            14'd16050: out = 14'h1055;
            14'd16051: out = 14'h1055;
            14'd16052: out = 14'h1055;
            14'd16053: out = 14'h1054;
            14'd16054: out = 14'h1054;
            14'd16055: out = 14'h1054;
            14'd16056: out = 14'h1054;
            14'd16057: out = 14'h1053;
            14'd16058: out = 14'h1053;
            14'd16059: out = 14'h1053;
            14'd16060: out = 14'h1053;
            14'd16061: out = 14'h1052;
            14'd16062: out = 14'h1052;
            14'd16063: out = 14'h1052;
            14'd16064: out = 14'h1052;
            14'd16065: out = 14'h1051;
            14'd16066: out = 14'h1051;
            14'd16067: out = 14'h1051;
            14'd16068: out = 14'h1051;
            14'd16069: out = 14'h1050;
            14'd16070: out = 14'h1050;
            14'd16071: out = 14'h1050;
            14'd16072: out = 14'h1050;
            14'd16073: out = 14'h104F;
            14'd16074: out = 14'h104F;
            14'd16075: out = 14'h104F;
            14'd16076: out = 14'h104E;
            14'd16077: out = 14'h104E;
            14'd16078: out = 14'h104E;
            14'd16079: out = 14'h104E;
            14'd16080: out = 14'h104D;
            14'd16081: out = 14'h104D;
            14'd16082: out = 14'h104D;
            14'd16083: out = 14'h104D;
            14'd16084: out = 14'h104C;
            14'd16085: out = 14'h104C;
            14'd16086: out = 14'h104C;
            14'd16087: out = 14'h104C;
            14'd16088: out = 14'h104B;
            14'd16089: out = 14'h104B;
            14'd16090: out = 14'h104B;
            14'd16091: out = 14'h104B;
            14'd16092: out = 14'h104A;
            14'd16093: out = 14'h104A;
            14'd16094: out = 14'h104A;
            14'd16095: out = 14'h104A;
            14'd16096: out = 14'h1049;
            14'd16097: out = 14'h1049;
            14'd16098: out = 14'h1049;
            14'd16099: out = 14'h1049;
            14'd16100: out = 14'h1048;
            14'd16101: out = 14'h1048;
            14'd16102: out = 14'h1048;
            14'd16103: out = 14'h1047;
            14'd16104: out = 14'h1047;
            14'd16105: out = 14'h1047;
            14'd16106: out = 14'h1047;
            14'd16107: out = 14'h1046;
            14'd16108: out = 14'h1046;
            14'd16109: out = 14'h1046;
            14'd16110: out = 14'h1046;
            14'd16111: out = 14'h1045;
            14'd16112: out = 14'h1045;
            14'd16113: out = 14'h1045;
            14'd16114: out = 14'h1045;
            14'd16115: out = 14'h1044;
            14'd16116: out = 14'h1044;
            14'd16117: out = 14'h1044;
            14'd16118: out = 14'h1044;
            14'd16119: out = 14'h1043;
            14'd16120: out = 14'h1043;
            14'd16121: out = 14'h1043;
            14'd16122: out = 14'h1043;
            14'd16123: out = 14'h1042;
            14'd16124: out = 14'h1042;
            14'd16125: out = 14'h1042;
            14'd16126: out = 14'h1042;
            14'd16127: out = 14'h1041;
            14'd16128: out = 14'h1041;
            14'd16129: out = 14'h1041;
            14'd16130: out = 14'h1040;
            14'd16131: out = 14'h1040;
            14'd16132: out = 14'h1040;
            14'd16133: out = 14'h1040;
            14'd16134: out = 14'h103F;
            14'd16135: out = 14'h103F;
            14'd16136: out = 14'h103F;
            14'd16137: out = 14'h103F;
            14'd16138: out = 14'h103E;
            14'd16139: out = 14'h103E;
            14'd16140: out = 14'h103E;
            14'd16141: out = 14'h103E;
            14'd16142: out = 14'h103D;
            14'd16143: out = 14'h103D;
            14'd16144: out = 14'h103D;
            14'd16145: out = 14'h103D;
            14'd16146: out = 14'h103C;
            14'd16147: out = 14'h103C;
            14'd16148: out = 14'h103C;
            14'd16149: out = 14'h103C;
            14'd16150: out = 14'h103B;
            14'd16151: out = 14'h103B;
            14'd16152: out = 14'h103B;
            14'd16153: out = 14'h103B;
            14'd16154: out = 14'h103A;
            14'd16155: out = 14'h103A;
            14'd16156: out = 14'h103A;
            14'd16157: out = 14'h103A;
            14'd16158: out = 14'h1039;
            14'd16159: out = 14'h1039;
            14'd16160: out = 14'h1039;
            14'd16161: out = 14'h1039;
            14'd16162: out = 14'h1038;
            14'd16163: out = 14'h1038;
            14'd16164: out = 14'h1038;
            14'd16165: out = 14'h1037;
            14'd16166: out = 14'h1037;
            14'd16167: out = 14'h1037;
            14'd16168: out = 14'h1037;
            14'd16169: out = 14'h1036;
            14'd16170: out = 14'h1036;
            14'd16171: out = 14'h1036;
            14'd16172: out = 14'h1036;
            14'd16173: out = 14'h1035;
            14'd16174: out = 14'h1035;
            14'd16175: out = 14'h1035;
            14'd16176: out = 14'h1035;
            14'd16177: out = 14'h1034;
            14'd16178: out = 14'h1034;
            14'd16179: out = 14'h1034;
            14'd16180: out = 14'h1034;
            14'd16181: out = 14'h1033;
            14'd16182: out = 14'h1033;
            14'd16183: out = 14'h1033;
            14'd16184: out = 14'h1033;
            14'd16185: out = 14'h1032;
            14'd16186: out = 14'h1032;
            14'd16187: out = 14'h1032;
            14'd16188: out = 14'h1032;
            14'd16189: out = 14'h1031;
            14'd16190: out = 14'h1031;
            14'd16191: out = 14'h1031;
            14'd16192: out = 14'h1031;
            14'd16193: out = 14'h1030;
            14'd16194: out = 14'h1030;
            14'd16195: out = 14'h1030;
            14'd16196: out = 14'h1030;
            14'd16197: out = 14'h102F;
            14'd16198: out = 14'h102F;
            14'd16199: out = 14'h102F;
            14'd16200: out = 14'h102F;
            14'd16201: out = 14'h102E;
            14'd16202: out = 14'h102E;
            14'd16203: out = 14'h102E;
            14'd16204: out = 14'h102D;
            14'd16205: out = 14'h102D;
            14'd16206: out = 14'h102D;
            14'd16207: out = 14'h102D;
            14'd16208: out = 14'h102C;
            14'd16209: out = 14'h102C;
            14'd16210: out = 14'h102C;
            14'd16211: out = 14'h102C;
            14'd16212: out = 14'h102B;
            14'd16213: out = 14'h102B;
            14'd16214: out = 14'h102B;
            14'd16215: out = 14'h102B;
            14'd16216: out = 14'h102A;
            14'd16217: out = 14'h102A;
            14'd16218: out = 14'h102A;
            14'd16219: out = 14'h102A;
            14'd16220: out = 14'h1029;
            14'd16221: out = 14'h1029;
            14'd16222: out = 14'h1029;
            14'd16223: out = 14'h1029;
            14'd16224: out = 14'h1028;
            14'd16225: out = 14'h1028;
            14'd16226: out = 14'h1028;
            14'd16227: out = 14'h1028;
            14'd16228: out = 14'h1027;
            14'd16229: out = 14'h1027;
            14'd16230: out = 14'h1027;
            14'd16231: out = 14'h1027;
            14'd16232: out = 14'h1026;
            14'd16233: out = 14'h1026;
            14'd16234: out = 14'h1026;
            14'd16235: out = 14'h1026;
            14'd16236: out = 14'h1025;
            14'd16237: out = 14'h1025;
            14'd16238: out = 14'h1025;
            14'd16239: out = 14'h1025;
            14'd16240: out = 14'h1024;
            14'd16241: out = 14'h1024;
            14'd16242: out = 14'h1024;
            14'd16243: out = 14'h1024;
            14'd16244: out = 14'h1023;
            14'd16245: out = 14'h1023;
            14'd16246: out = 14'h1023;
            14'd16247: out = 14'h1023;
            14'd16248: out = 14'h1022;
            14'd16249: out = 14'h1022;
            14'd16250: out = 14'h1022;
            14'd16251: out = 14'h1022;
            14'd16252: out = 14'h1021;
            14'd16253: out = 14'h1021;
            14'd16254: out = 14'h1021;
            14'd16255: out = 14'h1021;
            14'd16256: out = 14'h1020;
            14'd16257: out = 14'h1020;
            14'd16258: out = 14'h1020;
            14'd16259: out = 14'h101F;
            14'd16260: out = 14'h101F;
            14'd16261: out = 14'h101F;
            14'd16262: out = 14'h101F;
            14'd16263: out = 14'h101E;
            14'd16264: out = 14'h101E;
            14'd16265: out = 14'h101E;
            14'd16266: out = 14'h101E;
            14'd16267: out = 14'h101D;
            14'd16268: out = 14'h101D;
            14'd16269: out = 14'h101D;
            14'd16270: out = 14'h101D;
            14'd16271: out = 14'h101C;
            14'd16272: out = 14'h101C;
            14'd16273: out = 14'h101C;
            14'd16274: out = 14'h101C;
            14'd16275: out = 14'h101B;
            14'd16276: out = 14'h101B;
            14'd16277: out = 14'h101B;
            14'd16278: out = 14'h101B;
            14'd16279: out = 14'h101A;
            14'd16280: out = 14'h101A;
            14'd16281: out = 14'h101A;
            14'd16282: out = 14'h101A;
            14'd16283: out = 14'h1019;
            14'd16284: out = 14'h1019;
            14'd16285: out = 14'h1019;
            14'd16286: out = 14'h1019;
            14'd16287: out = 14'h1018;
            14'd16288: out = 14'h1018;
            14'd16289: out = 14'h1018;
            14'd16290: out = 14'h1018;
            14'd16291: out = 14'h1017;
            14'd16292: out = 14'h1017;
            14'd16293: out = 14'h1017;
            14'd16294: out = 14'h1017;
            14'd16295: out = 14'h1016;
            14'd16296: out = 14'h1016;
            14'd16297: out = 14'h1016;
            14'd16298: out = 14'h1016;
            14'd16299: out = 14'h1015;
            14'd16300: out = 14'h1015;
            14'd16301: out = 14'h1015;
            14'd16302: out = 14'h1015;
            14'd16303: out = 14'h1014;
            14'd16304: out = 14'h1014;
            14'd16305: out = 14'h1014;
            14'd16306: out = 14'h1014;
            14'd16307: out = 14'h1013;
            14'd16308: out = 14'h1013;
            14'd16309: out = 14'h1013;
            14'd16310: out = 14'h1013;
            14'd16311: out = 14'h1012;
            14'd16312: out = 14'h1012;
            14'd16313: out = 14'h1012;
            14'd16314: out = 14'h1012;
            14'd16315: out = 14'h1011;
            14'd16316: out = 14'h1011;
            14'd16317: out = 14'h1011;
            14'd16318: out = 14'h1011;
            14'd16319: out = 14'h1010;
            14'd16320: out = 14'h1010;
            14'd16321: out = 14'h1010;
            14'd16322: out = 14'h1010;
            14'd16323: out = 14'h100F;
            14'd16324: out = 14'h100F;
            14'd16325: out = 14'h100F;
            14'd16326: out = 14'h100F;
            14'd16327: out = 14'h100E;
            14'd16328: out = 14'h100E;
            14'd16329: out = 14'h100E;
            14'd16330: out = 14'h100E;
            14'd16331: out = 14'h100D;
            14'd16332: out = 14'h100D;
            14'd16333: out = 14'h100D;
            14'd16334: out = 14'h100D;
            14'd16335: out = 14'h100C;
            14'd16336: out = 14'h100C;
            14'd16337: out = 14'h100C;
            14'd16338: out = 14'h100C;
            14'd16339: out = 14'h100B;
            14'd16340: out = 14'h100B;
            14'd16341: out = 14'h100B;
            14'd16342: out = 14'h100B;
            14'd16343: out = 14'h100A;
            14'd16344: out = 14'h100A;
            14'd16345: out = 14'h100A;
            14'd16346: out = 14'h100A;
            14'd16347: out = 14'h1009;
            14'd16348: out = 14'h1009;
            14'd16349: out = 14'h1009;
            14'd16350: out = 14'h1009;
            14'd16351: out = 14'h1008;
            14'd16352: out = 14'h1008;
            14'd16353: out = 14'h1008;
            14'd16354: out = 14'h1008;
            14'd16355: out = 14'h1007;
            14'd16356: out = 14'h1007;
            14'd16357: out = 14'h1007;
            14'd16358: out = 14'h1007;
            14'd16359: out = 14'h1006;
            14'd16360: out = 14'h1006;
            14'd16361: out = 14'h1006;
            14'd16362: out = 14'h1006;
            14'd16363: out = 14'h1005;
            14'd16364: out = 14'h1005;
            14'd16365: out = 14'h1005;
            14'd16366: out = 14'h1005;
            14'd16367: out = 14'h1004;
            14'd16368: out = 14'h1004;
            14'd16369: out = 14'h1004;
            14'd16370: out = 14'h1004;
            14'd16371: out = 14'h1003;
            14'd16372: out = 14'h1003;
            14'd16373: out = 14'h1003;
            14'd16374: out = 14'h1003;
            14'd16375: out = 14'h1002;
            14'd16376: out = 14'h1002;
            14'd16377: out = 14'h1002;
            14'd16378: out = 14'h1002;
            14'd16379: out = 14'h1001;
            14'd16380: out = 14'h1001;
            14'd16381: out = 14'h1001;
            14'd16382: out = 14'h1001;
            14'd16383: out = 14'h1000;
            default: out = 14'h0000;
        endcase
        end
    end
endmodule
