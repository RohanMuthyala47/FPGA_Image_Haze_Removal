module Saturation_Correction_Multiplier (
    input  [15:0] x1,       // Ac^0.3 in Q8.8 format
    input  [15:0] x2,       // Jc^0.7 in Q8.8 format
    output [7:0]  result    // Final 8-bit saturation corrected pixel
);

    // Q8.8 * Q8.8 = Q16.16 result
    wire [31:0] mult_result = x1 * x2;

    // Extract the integer part from the Q16.16 fixed-point result
    assign result = mult_result[23:16];  // Scaling down to 8 bit value

endmodule
