module Atmospheric_Light_Reciprocal_LUT (
    input      [7:0] in,
    output reg [9:0] out
);

    always @(*) begin
        casez (in)
            8'd  1: out = 10'd1024;  // 1/1 ≈ 1.00000000
            8'd  2: out = 10'd 512;  // 1/2 ≈ 0.50000000
            8'd  3: out = 10'd 341;  // 1/3 ≈ 0.33333333
            8'd  4: out = 10'd 256;  // 1/4 ≈ 0.25000000
            8'd  5: out = 10'd 205;  // 1/5 ≈ 0.20000000
            8'd  6: out = 10'd 171;  // 1/6 ≈ 0.16666667
            8'd  7: out = 10'd 146;  // 1/7 ≈ 0.14285714
            8'd  8: out = 10'd 128;  // 1/8 ≈ 0.12500000
            8'd  9: out = 10'd 114;  // 1/9 ≈ 0.11111111
            8'd 10: out = 10'd 102;  // 1/10 ≈ 0.10000000
            8'd 11: out = 10'd  93;  // 1/11 ≈ 0.09090909
            8'd 12: out = 10'd  85;  // 1/12 ≈ 0.08333333
            8'd 13: out = 10'd  79;  // 1/13 ≈ 0.07692308
            8'd 14: out = 10'd  73;  // 1/14 ≈ 0.07142857
            8'd 15: out = 10'd  68;  // 1/15 ≈ 0.06666667
            8'd 16: out = 10'd  64;  // 1/16 ≈ 0.06250000
            8'd 17: out = 10'd  60;  // 1/17 ≈ 0.05882353
            8'd 18: out = 10'd  57;  // 1/18 ≈ 0.05555556
            8'd 19: out = 10'd  54;  // 1/19 ≈ 0.05263158
            8'd 20: out = 10'd  51;  // 1/20 ≈ 0.05000000
            8'd 21: out = 10'd  49;  // 1/21 ≈ 0.04761905
            8'd 22: out = 10'd  47;  // 1/22 ≈ 0.04545455
            8'd 23: out = 10'd  45;  // 1/23 ≈ 0.04347826
            8'd 24: out = 10'd  43;  // 1/24 ≈ 0.04166667
            8'd 25: out = 10'd  41;  // 1/25 ≈ 0.04000000
            8'd 26: out = 10'd  39;  // 1/26 ≈ 0.03846154
            8'd 27: out = 10'd  38;  // 1/27 ≈ 0.03703704
            8'd 28: out = 10'd  37;  // 1/28 ≈ 0.03571429
            8'd 29: out = 10'd  35;  // 1/29 ≈ 0.03448276
            8'd 30: out = 10'd  34;  // 1/30 ≈ 0.03333333
            8'd 31: out = 10'd  33;  // 1/31 ≈ 0.03225806
            8'd 32: out = 10'd  32;  // 1/32 ≈ 0.03125000
            8'd 33: out = 10'd  31;  // 1/33 ≈ 0.03030303
            8'd 34: out = 10'd  30;  // 1/34 ≈ 0.02941176
            8'd 35: out = 10'd  29;  // 1/35 ≈ 0.02857143
            8'd 36: out = 10'd  28;  // 1/36 ≈ 0.02777778
            8'd 37: out = 10'd  28;  // 1/37 ≈ 0.02702703
            8'd 38: out = 10'd  27;  // 1/38 ≈ 0.02631579
            8'd 39: out = 10'd  26;  // 1/39 ≈ 0.02564103
            8'd 40: out = 10'd  26;  // 1/40 ≈ 0.02500000
            8'd 41: out = 10'd  25;  // 1/41 ≈ 0.02439024
            8'd 42: out = 10'd  24;  // 1/42 ≈ 0.02380952
            8'd 43: out = 10'd  24;  // 1/43 ≈ 0.02325581
            8'd 44: out = 10'd  23;  // 1/44 ≈ 0.02272727
            8'd 45: out = 10'd  23;  // 1/45 ≈ 0.02222222
            8'd 46: out = 10'd  22;  // 1/46 ≈ 0.02173913
            8'd 47: out = 10'd  22;  // 1/47 ≈ 0.02127660
            8'd 48: out = 10'd  21;  // 1/48 ≈ 0.02083333
            8'd 49: out = 10'd  21;  // 1/49 ≈ 0.02040816
            8'd 50: out = 10'd  20;  // 1/50 ≈ 0.02000000
            8'd 51: out = 10'd  20;  // 1/51 ≈ 0.01960784
            8'd 52: out = 10'd  20;  // 1/52 ≈ 0.01923077
            8'd 53: out = 10'd  19;  // 1/53 ≈ 0.01886792
            8'd 54: out = 10'd  19;  // 1/54 ≈ 0.01851852
            8'd 55: out = 10'd  19;  // 1/55 ≈ 0.01818182
            8'd 56: out = 10'd  18;  // 1/56 ≈ 0.01785714
            8'd 57: out = 10'd  18;  // 1/57 ≈ 0.01754386
            8'd 58: out = 10'd  18;  // 1/58 ≈ 0.01724138
            8'd 59: out = 10'd  17;  // 1/59 ≈ 0.01694915
            8'd 60: out = 10'd  17;  // 1/60 ≈ 0.01666667
            8'd 61: out = 10'd  17;  // 1/61 ≈ 0.01639344
            8'd 62: out = 10'd  17;  // 1/62 ≈ 0.01612903
            8'd 63: out = 10'd  16;  // 1/63 ≈ 0.01587302
            8'd 64: out = 10'd  16;  // 1/64 ≈ 0.01562500
            8'd 65: out = 10'd  16;  // 1/65 ≈ 0.01538462
            8'd 66: out = 10'd  16;  // 1/66 ≈ 0.01515152
            8'd 67: out = 10'd  15;  // 1/67 ≈ 0.01492537
            8'd 68: out = 10'd  15;  // 1/68 ≈ 0.01470588
            8'd 69: out = 10'd  15;  // 1/69 ≈ 0.01449275
            8'd 70: out = 10'd  15;  // 1/70 ≈ 0.01428571
            8'd 71: out = 10'd  14;  // 1/71 ≈ 0.01408451
            8'd 72: out = 10'd  14;  // 1/72 ≈ 0.01388889
            8'd 73: out = 10'd  14;  // 1/73 ≈ 0.01369863
            8'd 74: out = 10'd  14;  // 1/74 ≈ 0.01351351
            8'd 75: out = 10'd  14;  // 1/75 ≈ 0.01333333
            8'd 76: out = 10'd  13;  // 1/76 ≈ 0.01315789
            8'd 77: out = 10'd  13;  // 1/77 ≈ 0.01298701
            8'd 78: out = 10'd  13;  // 1/78 ≈ 0.01282051
            8'd 79: out = 10'd  13;  // 1/79 ≈ 0.01265823
            8'd 80: out = 10'd  13;  // 1/80 ≈ 0.01250000
            8'd 81: out = 10'd  13;  // 1/81 ≈ 0.01234568
            8'd 82: out = 10'd  12;  // 1/82 ≈ 0.01219512
            8'd 83: out = 10'd  12;  // 1/83 ≈ 0.01204819
            8'd 84: out = 10'd  12;  // 1/84 ≈ 0.01190476
            8'd 85: out = 10'd  12;  // 1/85 ≈ 0.01176471
            8'd 86: out = 10'd  12;  // 1/86 ≈ 0.01162791
            8'd 87: out = 10'd  12;  // 1/87 ≈ 0.01149425
            8'd 88: out = 10'd  12;  // 1/88 ≈ 0.01136364
            8'd 89: out = 10'd  12;  // 1/89 ≈ 0.01123596
            8'd 90: out = 10'd  11;  // 1/90 ≈ 0.01111111
            8'd 91: out = 10'd  11;  // 1/91 ≈ 0.01098901
            8'd 92: out = 10'd  11;  // 1/92 ≈ 0.01086957
            8'd 93: out = 10'd  11;  // 1/93 ≈ 0.01075269
            8'd 94: out = 10'd  11;  // 1/94 ≈ 0.01063830
            8'd 95: out = 10'd  11;  // 1/95 ≈ 0.01052632
            8'd 96: out = 10'd  11;  // 1/96 ≈ 0.01041667
            8'd 97: out = 10'd  11;  // 1/97 ≈ 0.01030928
            8'd 98: out = 10'd  10;  // 1/98 ≈ 0.01020408
            8'd 99: out = 10'd  10;  // 1/99 ≈ 0.01010101
            8'd100: out = 10'd  10;  // 1/100 ≈ 0.01000000
            8'd101: out = 10'd  10;  // 1/101 ≈ 0.00990099
            8'd102: out = 10'd  10;  // 1/102 ≈ 0.00980392
            8'd103: out = 10'd  10;  // 1/103 ≈ 0.00970874
            8'd104: out = 10'd  10;  // 1/104 ≈ 0.00961538
            8'd105: out = 10'd  10;  // 1/105 ≈ 0.00952381
            8'd106: out = 10'd  10;  // 1/106 ≈ 0.00943396
            8'd107: out = 10'd  10;  // 1/107 ≈ 0.00934579
            8'd108: out = 10'd   9;  // 1/108 ≈ 0.00925926
            8'd109: out = 10'd   9;  // 1/109 ≈ 0.00917431
            8'd110: out = 10'd   9;  // 1/110 ≈ 0.00909091
            8'd111: out = 10'd   9;  // 1/111 ≈ 0.00900901
            8'd112: out = 10'd   9;  // 1/112 ≈ 0.00892857
            8'd113: out = 10'd   9;  // 1/113 ≈ 0.00884956
            8'd114: out = 10'd   9;  // 1/114 ≈ 0.00877193
            8'd115: out = 10'd   9;  // 1/115 ≈ 0.00869565
            8'd116: out = 10'd   9;  // 1/116 ≈ 0.00862069
            8'd117: out = 10'd   9;  // 1/117 ≈ 0.00854701
            8'd118: out = 10'd   9;  // 1/118 ≈ 0.00847458
            8'd119: out = 10'd   9;  // 1/119 ≈ 0.00840336
            8'd120: out = 10'd   9;  // 1/120 ≈ 0.00833333
            8'd121: out = 10'd   8;  // 1/121 ≈ 0.00826446
            8'd122: out = 10'd   8;  // 1/122 ≈ 0.00819672
            8'd123: out = 10'd   8;  // 1/123 ≈ 0.00813008
            8'd124: out = 10'd   8;  // 1/124 ≈ 0.00806452
            8'd125: out = 10'd   8;  // 1/125 ≈ 0.00800000
            8'd126: out = 10'd   8;  // 1/126 ≈ 0.00793651
            8'd127: out = 10'd   8;  // 1/127 ≈ 0.00787402
            8'd128: out = 10'd   8;  // 1/128 ≈ 0.00781250
            8'd129: out = 10'd   8;  // 1/129 ≈ 0.00775194
            8'd130: out = 10'd   8;  // 1/130 ≈ 0.00769231
            8'd131: out = 10'd   8;  // 1/131 ≈ 0.00763359
            8'd132: out = 10'd   8;  // 1/132 ≈ 0.00757576
            8'd133: out = 10'd   8;  // 1/133 ≈ 0.00751880
            8'd134: out = 10'd   8;  // 1/134 ≈ 0.00746269
            8'd135: out = 10'd   8;  // 1/135 ≈ 0.00740741
            8'd136: out = 10'd   8;  // 1/136 ≈ 0.00735294
            8'd137: out = 10'd   7;  // 1/137 ≈ 0.00729927
            8'd138: out = 10'd   7;  // 1/138 ≈ 0.00724638
            8'd139: out = 10'd   7;  // 1/139 ≈ 0.00719424
            8'd140: out = 10'd   7;  // 1/140 ≈ 0.00714286
            8'd141: out = 10'd   7;  // 1/141 ≈ 0.00709220
            8'd142: out = 10'd   7;  // 1/142 ≈ 0.00704225
            8'd143: out = 10'd   7;  // 1/143 ≈ 0.00699301
            8'd144: out = 10'd   7;  // 1/144 ≈ 0.00694444
            8'd145: out = 10'd   7;  // 1/145 ≈ 0.00689655
            8'd146: out = 10'd   7;  // 1/146 ≈ 0.00684932
            8'd147: out = 10'd   7;  // 1/147 ≈ 0.00680272
            8'd148: out = 10'd   7;  // 1/148 ≈ 0.00675676
            8'd149: out = 10'd   7;  // 1/149 ≈ 0.00671141
            8'd150: out = 10'd   7;  // 1/150 ≈ 0.00666667
            8'd151: out = 10'd   7;  // 1/151 ≈ 0.00662252
            8'd152: out = 10'd   7;  // 1/152 ≈ 0.00657895
            8'd153: out = 10'd   7;  // 1/153 ≈ 0.00653595
            8'd154: out = 10'd   7;  // 1/154 ≈ 0.00649351
            8'd155: out = 10'd   7;  // 1/155 ≈ 0.00645161
            8'd156: out = 10'd   7;  // 1/156 ≈ 0.00641026
            8'd157: out = 10'd   7;  // 1/157 ≈ 0.00636943
            8'd158: out = 10'd   6;  // 1/158 ≈ 0.00632911
            8'd159: out = 10'd   6;  // 1/159 ≈ 0.00628931
            8'd160: out = 10'd   6;  // 1/160 ≈ 0.00625000
            8'd161: out = 10'd   6;  // 1/161 ≈ 0.00621118
            8'd162: out = 10'd   6;  // 1/162 ≈ 0.00617284
            8'd163: out = 10'd   6;  // 1/163 ≈ 0.00613497
            8'd164: out = 10'd   6;  // 1/164 ≈ 0.00609756
            8'd165: out = 10'd   6;  // 1/165 ≈ 0.00606061
            8'd166: out = 10'd   6;  // 1/166 ≈ 0.00602410
            8'd167: out = 10'd   6;  // 1/167 ≈ 0.00598802
            8'd168: out = 10'd   6;  // 1/168 ≈ 0.00595238
            8'd169: out = 10'd   6;  // 1/169 ≈ 0.00591716
            8'd170: out = 10'd   6;  // 1/170 ≈ 0.00588235
            8'd171: out = 10'd   6;  // 1/171 ≈ 0.00584795
            8'd172: out = 10'd   6;  // 1/172 ≈ 0.00581395
            8'd173: out = 10'd   6;  // 1/173 ≈ 0.00578035
            8'd174: out = 10'd   6;  // 1/174 ≈ 0.00574713
            8'd175: out = 10'd   6;  // 1/175 ≈ 0.00571429
            8'd176: out = 10'd   6;  // 1/176 ≈ 0.00568182
            8'd177: out = 10'd   6;  // 1/177 ≈ 0.00564972
            8'd178: out = 10'd   6;  // 1/178 ≈ 0.00561798
            8'd179: out = 10'd   6;  // 1/179 ≈ 0.00558659
            8'd180: out = 10'd   6;  // 1/180 ≈ 0.00555556
            8'd181: out = 10'd   6;  // 1/181 ≈ 0.00552486
            8'd182: out = 10'd   6;  // 1/182 ≈ 0.00549451
            8'd183: out = 10'd   6;  // 1/183 ≈ 0.00546448
            8'd184: out = 10'd   6;  // 1/184 ≈ 0.00543478
            8'd185: out = 10'd   6;  // 1/185 ≈ 0.00540541
            8'd186: out = 10'd   6;  // 1/186 ≈ 0.00537634
            8'd187: out = 10'd   5;  // 1/187 ≈ 0.00534759
            8'd188: out = 10'd   5;  // 1/188 ≈ 0.00531915
            8'd189: out = 10'd   5;  // 1/189 ≈ 0.00529101
            8'd190: out = 10'd   5;  // 1/190 ≈ 0.00526316
            8'd191: out = 10'd   5;  // 1/191 ≈ 0.00523560
            8'd192: out = 10'd   5;  // 1/192 ≈ 0.00520833
            8'd193: out = 10'd   5;  // 1/193 ≈ 0.00518135
            8'd194: out = 10'd   5;  // 1/194 ≈ 0.00515464
            8'd195: out = 10'd   5;  // 1/195 ≈ 0.00512821
            8'd196: out = 10'd   5;  // 1/196 ≈ 0.00510204
            8'd197: out = 10'd   5;  // 1/197 ≈ 0.00507614
            8'd198: out = 10'd   5;  // 1/198 ≈ 0.00505051
            8'd199: out = 10'd   5;  // 1/199 ≈ 0.00502513
            8'd200: out = 10'd   5;  // 1/200 ≈ 0.00500000
            8'd201: out = 10'd   5;  // 1/201 ≈ 0.00497512
            8'd202: out = 10'd   5;  // 1/202 ≈ 0.00495050
            8'd203: out = 10'd   5;  // 1/203 ≈ 0.00492611
            8'd204: out = 10'd   5;  // 1/204 ≈ 0.00490196
            8'd205: out = 10'd   5;  // 1/205 ≈ 0.00487805
            8'd206: out = 10'd   5;  // 1/206 ≈ 0.00485437
            8'd207: out = 10'd   5;  // 1/207 ≈ 0.00483092
            8'd208: out = 10'd   5;  // 1/208 ≈ 0.00480769
            8'd209: out = 10'd   5;  // 1/209 ≈ 0.00478469
            8'd210: out = 10'd   5;  // 1/210 ≈ 0.00476190
            8'd211: out = 10'd   5;  // 1/211 ≈ 0.00473934
            8'd212: out = 10'd   5;  // 1/212 ≈ 0.00471698
            8'd213: out = 10'd   5;  // 1/213 ≈ 0.00469484
            8'd214: out = 10'd   5;  // 1/214 ≈ 0.00467290
            8'd215: out = 10'd   5;  // 1/215 ≈ 0.00465116
            8'd216: out = 10'd   5;  // 1/216 ≈ 0.00462963
            8'd217: out = 10'd   5;  // 1/217 ≈ 0.00460829
            8'd218: out = 10'd   5;  // 1/218 ≈ 0.00458716
            8'd219: out = 10'd   5;  // 1/219 ≈ 0.00456621
            8'd220: out = 10'd   5;  // 1/220 ≈ 0.00454545
            8'd221: out = 10'd   5;  // 1/221 ≈ 0.00452489
            8'd222: out = 10'd   5;  // 1/222 ≈ 0.00450450
            8'd223: out = 10'd   5;  // 1/223 ≈ 0.00448430
            8'd224: out = 10'd   5;  // 1/224 ≈ 0.00446429
            8'd225: out = 10'd   5;  // 1/225 ≈ 0.00444444
            8'd226: out = 10'd   5;  // 1/226 ≈ 0.00442478
            8'd227: out = 10'd   5;  // 1/227 ≈ 0.00440529
            8'd228: out = 10'd   4;  // 1/228 ≈ 0.00438596
            8'd229: out = 10'd   4;  // 1/229 ≈ 0.00436681
            8'd230: out = 10'd   4;  // 1/230 ≈ 0.00434783
            8'd231: out = 10'd   4;  // 1/231 ≈ 0.00432900
            8'd232: out = 10'd   4;  // 1/232 ≈ 0.00431034
            8'd233: out = 10'd   4;  // 1/233 ≈ 0.00429185
            8'd234: out = 10'd   4;  // 1/234 ≈ 0.00427350
            8'd235: out = 10'd   4;  // 1/235 ≈ 0.00425532
            8'd236: out = 10'd   4;  // 1/236 ≈ 0.00423729
            8'd237: out = 10'd   4;  // 1/237 ≈ 0.00421941
            8'd238: out = 10'd   4;  // 1/238 ≈ 0.00420168
            8'd239: out = 10'd   4;  // 1/239 ≈ 0.00418410
            8'd240: out = 10'd   4;  // 1/240 ≈ 0.00416667
            8'd241: out = 10'd   4;  // 1/241 ≈ 0.00414938
            8'd242: out = 10'd   4;  // 1/242 ≈ 0.00413223
            8'd243: out = 10'd   4;  // 1/243 ≈ 0.00411523
            8'd244: out = 10'd   4;  // 1/244 ≈ 0.00409836
            8'd245: out = 10'd   4;  // 1/245 ≈ 0.00408163
            8'd246: out = 10'd   4;  // 1/246 ≈ 0.00406504
            8'd247: out = 10'd   4;  // 1/247 ≈ 0.00404858
            8'd248: out = 10'd   4;  // 1/248 ≈ 0.00403226
            8'd249: out = 10'd   4;  // 1/249 ≈ 0.00401606
            8'd250: out = 10'd   4;  // 1/250 ≈ 0.00400000
            8'd251: out = 10'd   4;  // 1/251 ≈ 0.00398406
            8'd252: out = 10'd   4;  // 1/252 ≈ 0.00396825
            8'd253: out = 10'd   4;  // 1/253 ≈ 0.00395257
            8'd254: out = 10'd   4;  // 1/254 ≈ 0.00393701
            8'd255: out = 10'd   4;  // 1/255 ≈ 0.00392157
            default: out = 10'd1023; // undefined for 0
        endcase
    end

endmodule
