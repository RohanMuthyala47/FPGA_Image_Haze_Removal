// Look Up Tables for applying saturation correction

// LUT for x^0.35 in Q3.9 format
module LUT_035 (
    input      [7:0] in,  // Q8.0 input
    output reg [11:0] out // Q3.9 output
);

    always @(*) begin
        case (in)
            8'd0  : out = 12'd0;  // 0^0.35 ~= 0.000000
            8'd1  : out = 12'd512;  // 1^0.35 ~= 1.000000
            8'd2  : out = 12'd653;  // 2^0.35 ~= 1.274561
            8'd3  : out = 12'd752;  // 3^0.35 ~= 1.468901
            8'd4  : out = 12'd832;  // 4^0.35 ~= 1.624505
            8'd5  : out = 12'd899;  // 5^0.35 ~= 1.756465
            8'd6  : out = 12'd959;  // 6^0.35 ~= 1.872203
            8'd7  : out = 12'd1012;  // 7^0.35 ~= 1.975988
            8'd8  : out = 12'd1060;  // 8^0.35 ~= 2.070530
            8'd9  : out = 12'd1105;  // 9^0.35 ~= 2.157669
            8'd10 : out = 12'd1146;  // 10^0.35 ~= 2.238721
            8'd11 : out = 12'd1185;  // 11^0.35 ~= 2.314661
            8'd12 : out = 12'd1222;  // 12^0.35 ~= 2.386236
            8'd13 : out = 12'd1256;  // 13^0.35 ~= 2.454032
            8'd14 : out = 12'd1289;  // 14^0.35 ~= 2.518517
            8'd15 : out = 12'd1321;  // 15^0.35 ~= 2.580073
            8'd16 : out = 12'd1351;  // 16^0.35 ~= 2.639016
            8'd17 : out = 12'd1380;  // 17^0.35 ~= 2.695610
            8'd18 : out = 12'd1408;  // 18^0.35 ~= 2.750080
            8'd19 : out = 12'd1435;  // 19^0.35 ~= 2.802617
            8'd20 : out = 12'd1461;  // 20^0.35 ~= 2.853386
            8'd21 : out = 12'd1486;  // 21^0.35 ~= 2.902530
            8'd22 : out = 12'd1510;  // 22^0.35 ~= 2.950176
            8'd23 : out = 12'd1534;  // 23^0.35 ~= 2.996434
            8'd24 : out = 12'd1557;  // 24^0.35 ~= 3.041403
            8'd25 : out = 12'd1580;  // 25^0.35 ~= 3.085169
            8'd26 : out = 12'd1601;  // 26^0.35 ~= 3.127812
            8'd27 : out = 12'd1623;  // 27^0.35 ~= 3.169402
            8'd28 : out = 12'd1644;  // 28^0.35 ~= 3.210002
            8'd29 : out = 12'd1664;  // 29^0.35 ~= 3.249670
            8'd30 : out = 12'd1684;  // 30^0.35 ~= 3.288459
            8'd31 : out = 12'd1703;  // 31^0.35 ~= 3.326416
            8'd32 : out = 12'd1722;  // 32^0.35 ~= 3.363586
            8'd33 : out = 12'd1741;  // 33^0.35 ~= 3.400008
            8'd34 : out = 12'd1759;  // 34^0.35 ~= 3.435719
            8'd35 : out = 12'd1777;  // 35^0.35 ~= 3.470754
            8'd36 : out = 12'd1795;  // 36^0.35 ~= 3.505144
            8'd37 : out = 12'd1812;  // 37^0.35 ~= 3.538919
            8'd38 : out = 12'd1829;  // 38^0.35 ~= 3.572105
            8'd39 : out = 12'd1846;  // 39^0.35 ~= 3.604729
            8'd40 : out = 12'd1862;  // 40^0.35 ~= 3.636813
            8'd41 : out = 12'd1878;  // 41^0.35 ~= 3.668380
            8'd42 : out = 12'd1894;  // 42^0.35 ~= 3.699451
            8'd43 : out = 12'd1910;  // 43^0.35 ~= 3.730044
            8'd44 : out = 12'd1925;  // 44^0.35 ~= 3.760178
            8'd45 : out = 12'd1940;  // 45^0.35 ~= 3.789871
            8'd46 : out = 12'd1955;  // 46^0.35 ~= 3.819137
            8'd47 : out = 12'd1970;  // 47^0.35 ~= 3.847993
            8'd48 : out = 12'd1985;  // 48^0.35 ~= 3.876452
            8'd49 : out = 12'd1999;  // 49^0.35 ~= 3.904529
            8'd50 : out = 12'd2013;  // 50^0.35 ~= 3.932235
            8'd51 : out = 12'd2027;  // 51^0.35 ~= 3.959584
            8'd52 : out = 12'd2041;  // 52^0.35 ~= 3.986586
            8'd53 : out = 12'd2055;  // 53^0.35 ~= 4.013253
            8'd54 : out = 12'd2068;  // 54^0.35 ~= 4.039595
            8'd55 : out = 12'd2082;  // 55^0.35 ~= 4.065621
            8'd56 : out = 12'd2095;  // 56^0.35 ~= 4.091342
            8'd57 : out = 12'd2108;  // 57^0.35 ~= 4.116766
            8'd58 : out = 12'd2121;  // 58^0.35 ~= 4.141902
            8'd59 : out = 12'd2133;  // 59^0.35 ~= 4.166757
            8'd60 : out = 12'd2146;  // 60^0.35 ~= 4.191340
            8'd61 : out = 12'd2158;  // 61^0.35 ~= 4.215659
            8'd62 : out = 12'd2171;  // 62^0.35 ~= 4.239719
            8'd63 : out = 12'd2183;  // 63^0.35 ~= 4.263529
            8'd64 : out = 12'd2195;  // 64^0.35 ~= 4.287094
            8'd65 : out = 12'd2207;  // 65^0.35 ~= 4.310421
            8'd66 : out = 12'd2219;  // 66^0.35 ~= 4.333516
            8'd67 : out = 12'd2230;  // 67^0.35 ~= 4.356384
            8'd68 : out = 12'd2242;  // 68^0.35 ~= 4.379032
            8'd69 : out = 12'd2254;  // 69^0.35 ~= 4.401464
            8'd70 : out = 12'd2265;  // 70^0.35 ~= 4.423686
            8'd71 : out = 12'd2276;  // 71^0.35 ~= 4.445703
            8'd72 : out = 12'd2287;  // 72^0.35 ~= 4.467519
            8'd73 : out = 12'd2298;  // 73^0.35 ~= 4.489138
            8'd74 : out = 12'd2309;  // 74^0.35 ~= 4.510567
            8'd75 : out = 12'd2320;  // 75^0.35 ~= 4.531807
            8'd76 : out = 12'd2331;  // 76^0.35 ~= 4.552865
            8'd77 : out = 12'd2342;  // 77^0.35 ~= 4.573743
            8'd78 : out = 12'd2352;  // 78^0.35 ~= 4.594446
            8'd79 : out = 12'd2363;  // 79^0.35 ~= 4.614976
            8'd80 : out = 12'd2373;  // 80^0.35 ~= 4.635339
            8'd81 : out = 12'd2384;  // 81^0.35 ~= 4.655537
            8'd82 : out = 12'd2394;  // 82^0.35 ~= 4.675573
            8'd83 : out = 12'd2404;  // 83^0.35 ~= 4.695451
            8'd84 : out = 12'd2414;  // 84^0.35 ~= 4.715174
            8'd85 : out = 12'd2424;  // 85^0.35 ~= 4.734745
            8'd86 : out = 12'd2434;  // 86^0.35 ~= 4.754167
            8'd87 : out = 12'd2444;  // 87^0.35 ~= 4.773443
            8'd88 : out = 12'd2454;  // 88^0.35 ~= 4.792575
            8'd89 : out = 12'd2464;  // 89^0.35 ~= 4.811567
            8'd90 : out = 12'd2473;  // 90^0.35 ~= 4.830420
            8'd91 : out = 12'd2483;  // 91^0.35 ~= 4.849137
            8'd92 : out = 12'd2492;  // 92^0.35 ~= 4.867722
            8'd93 : out = 12'd2502;  // 93^0.35 ~= 4.886175
            8'd94 : out = 12'd2511;  // 94^0.35 ~= 4.904500
            8'd95 : out = 12'd2520;  // 95^0.35 ~= 4.922699
            8'd96 : out = 12'd2530;  // 96^0.35 ~= 4.940773
            8'd97 : out = 12'd2539;  // 97^0.35 ~= 4.958726
            8'd98 : out = 12'd2548;  // 98^0.35 ~= 4.976559
            8'd99 : out = 12'd2557;  // 99^0.35 ~= 4.994273
            8'd100: out = 12'd2566;  // 100^0.35 ~= 5.011872
            8'd101: out = 12'd2575;  // 101^0.35 ~= 5.029357
            8'd102: out = 12'd2584;  // 102^0.35 ~= 5.046730
            8'd103: out = 12'd2593;  // 103^0.35 ~= 5.063992
            8'd104: out = 12'd2602;  // 104^0.35 ~= 5.081146
            8'd105: out = 12'd2610;  // 105^0.35 ~= 5.098193
            8'd106: out = 12'd2619;  // 106^0.35 ~= 5.115134
            8'd107: out = 12'd2628;  // 107^0.35 ~= 5.131973
            8'd108: out = 12'd2636;  // 108^0.35 ~= 5.148709
            8'd109: out = 12'd2645;  // 109^0.35 ~= 5.165344
            8'd110: out = 12'd2653;  // 110^0.35 ~= 5.181881
            8'd111: out = 12'd2662;  // 111^0.35 ~= 5.198320
            8'd112: out = 12'd2670;  // 112^0.35 ~= 5.214664
            8'd113: out = 12'd2678;  // 113^0.35 ~= 5.230912
            8'd114: out = 12'd2686;  // 114^0.35 ~= 5.247068
            8'd115: out = 12'd2695;  // 115^0.35 ~= 5.263132
            8'd116: out = 12'd2703;  // 116^0.35 ~= 5.279105
            8'd117: out = 12'd2711;  // 117^0.35 ~= 5.294989
            8'd118: out = 12'd2719;  // 118^0.35 ~= 5.310785
            8'd119: out = 12'd2727;  // 119^0.35 ~= 5.326494
            8'd120: out = 12'd2735;  // 120^0.35 ~= 5.342118
            8'd121: out = 12'd2743;  // 121^0.35 ~= 5.357657
            8'd122: out = 12'd2751;  // 122^0.35 ~= 5.373113
            8'd123: out = 12'd2759;  // 123^0.35 ~= 5.388486
            8'd124: out = 12'd2767;  // 124^0.35 ~= 5.403779
            8'd125: out = 12'd2775;  // 125^0.35 ~= 5.418992
            8'd126: out = 12'd2782;  // 126^0.35 ~= 5.434126
            8'd127: out = 12'd2790;  // 127^0.35 ~= 5.449182
            8'd128: out = 12'd2798;  // 128^0.35 ~= 5.464161
            8'd129: out = 12'd2805;  // 129^0.35 ~= 5.479064
            8'd130: out = 12'd2813;  // 130^0.35 ~= 5.493893
            8'd131: out = 12'd2820;  // 131^0.35 ~= 5.508647
            8'd132: out = 12'd2828;  // 132^0.35 ~= 5.523329
            8'd133: out = 12'd2835;  // 133^0.35 ~= 5.537938
            8'd134: out = 12'd2843;  // 134^0.35 ~= 5.552476
            8'd135: out = 12'd2850;  // 135^0.35 ~= 5.566944
            8'd136: out = 12'd2858;  // 136^0.35 ~= 5.581342
            8'd137: out = 12'd2865;  // 137^0.35 ~= 5.595671
            8'd138: out = 12'd2872;  // 138^0.35 ~= 5.609933
            8'd139: out = 12'd2880;  // 139^0.35 ~= 5.624128
            8'd140: out = 12'd2887;  // 140^0.35 ~= 5.638256
            8'd141: out = 12'd2894;  // 141^0.35 ~= 5.652319
            8'd142: out = 12'd2901;  // 142^0.35 ~= 5.666318
            8'd143: out = 12'd2908;  // 143^0.35 ~= 5.680252
            8'd144: out = 12'd2915;  // 144^0.35 ~= 5.694123
            8'd145: out = 12'd2922;  // 145^0.35 ~= 5.707932
            8'd146: out = 12'd2929;  // 146^0.35 ~= 5.721679
            8'd147: out = 12'd2937;  // 147^0.35 ~= 5.735365
            8'd148: out = 12'd2943;  // 148^0.35 ~= 5.748991
            8'd149: out = 12'd2950;  // 149^0.35 ~= 5.762556
            8'd150: out = 12'd2957;  // 150^0.35 ~= 5.776063
            8'd151: out = 12'd2964;  // 151^0.35 ~= 5.789512
            8'd152: out = 12'd2971;  // 152^0.35 ~= 5.802902
            8'd153: out = 12'd2978;  // 153^0.35 ~= 5.816236
            8'd154: out = 12'd2985;  // 154^0.35 ~= 5.829513
            8'd155: out = 12'd2991;  // 155^0.35 ~= 5.842734
            8'd156: out = 12'd2998;  // 156^0.35 ~= 5.855899
            8'd157: out = 12'd3005;  // 157^0.35 ~= 5.869010
            8'd158: out = 12'd3012;  // 158^0.35 ~= 5.882067
            8'd159: out = 12'd3018;  // 159^0.35 ~= 5.895070
            8'd160: out = 12'd3025;  // 160^0.35 ~= 5.908021
            8'd161: out = 12'd3032;  // 161^0.35 ~= 5.920918
            8'd162: out = 12'd3038;  // 162^0.35 ~= 5.933764
            8'd163: out = 12'd3045;  // 163^0.35 ~= 5.946558
            8'd164: out = 12'd3051;  // 164^0.35 ~= 5.959301
            8'd165: out = 12'd3058;  // 165^0.35 ~= 5.971994
            8'd166: out = 12'd3064;  // 166^0.35 ~= 5.984637
            8'd167: out = 12'd3071;  // 167^0.35 ~= 5.997231
            8'd168: out = 12'd3077;  // 168^0.35 ~= 6.009775
            8'd169: out = 12'd3083;  // 169^0.35 ~= 6.022272
            8'd170: out = 12'd3090;  // 170^0.35 ~= 6.034720
            8'd171: out = 12'd3096;  // 171^0.35 ~= 6.047121
            8'd172: out = 12'd3102;  // 172^0.35 ~= 6.059474
            8'd173: out = 12'd3109;  // 173^0.35 ~= 6.071782
            8'd174: out = 12'd3115;  // 174^0.35 ~= 6.084042
            8'd175: out = 12'd3121;  // 175^0.35 ~= 6.096258
            8'd176: out = 12'd3128;  // 176^0.35 ~= 6.108428
            8'd177: out = 12'd3134;  // 177^0.35 ~= 6.120553
            8'd178: out = 12'd3140;  // 178^0.35 ~= 6.132633
            8'd179: out = 12'd3146;  // 179^0.35 ~= 6.144670
            8'd180: out = 12'd3152;  // 180^0.35 ~= 6.156663
            8'd181: out = 12'd3158;  // 181^0.35 ~= 6.168613
            8'd182: out = 12'd3164;  // 182^0.35 ~= 6.180520
            8'd183: out = 12'd3171;  // 183^0.35 ~= 6.192384
            8'd184: out = 12'd3177;  // 184^0.35 ~= 6.204206
            8'd185: out = 12'd3183;  // 185^0.35 ~= 6.215987
            8'd186: out = 12'd3189;  // 186^0.35 ~= 6.227726
            8'd187: out = 12'd3195;  // 187^0.35 ~= 6.239425
            8'd188: out = 12'd3201;  // 188^0.35 ~= 6.251083
            8'd189: out = 12'd3207;  // 189^0.35 ~= 6.262700
            8'd190: out = 12'd3212;  // 190^0.35 ~= 6.274278
            8'd191: out = 12'd3218;  // 191^0.35 ~= 6.285816
            8'd192: out = 12'd3224;  // 192^0.35 ~= 6.297315
            8'd193: out = 12'd3230;  // 193^0.35 ~= 6.308775
            8'd194: out = 12'd3236;  // 194^0.35 ~= 6.320197
            8'd195: out = 12'd3242;  // 195^0.35 ~= 6.331580
            8'd196: out = 12'd3248;  // 196^0.35 ~= 6.342926
            8'd197: out = 12'd3253;  // 197^0.35 ~= 6.354234
            8'd198: out = 12'd3259;  // 198^0.35 ~= 6.365504
            8'd199: out = 12'd3265;  // 199^0.35 ~= 6.376738
            8'd200: out = 12'd3271;  // 200^0.35 ~= 6.387935
            8'd201: out = 12'd3276;  // 201^0.35 ~= 6.399096
            8'd202: out = 12'd3282;  // 202^0.35 ~= 6.410221
            8'd203: out = 12'd3288;  // 203^0.35 ~= 6.421310
            8'd204: out = 12'd3293;  // 204^0.35 ~= 6.432363
            8'd205: out = 12'd3299;  // 205^0.35 ~= 6.443382
            8'd206: out = 12'd3305;  // 206^0.35 ~= 6.454365
            8'd207: out = 12'd3310;  // 207^0.35 ~= 6.465314
            8'd208: out = 12'd3316;  // 208^0.35 ~= 6.476229
            8'd209: out = 12'd3321;  // 209^0.35 ~= 6.487109
            8'd210: out = 12'd3327;  // 210^0.35 ~= 6.497956
            8'd211: out = 12'd3332;  // 211^0.35 ~= 6.508769
            8'd212: out = 12'd3338;  // 212^0.35 ~= 6.519549
            8'd213: out = 12'd3344;  // 213^0.35 ~= 6.530296
            8'd214: out = 12'd3349;  // 214^0.35 ~= 6.541010
            8'd215: out = 12'd3354;  // 215^0.35 ~= 6.551692
            8'd216: out = 12'd3360;  // 216^0.35 ~= 6.562341
            8'd217: out = 12'd3365;  // 217^0.35 ~= 6.572959
            8'd218: out = 12'd3371;  // 218^0.35 ~= 6.583544
            8'd219: out = 12'd3376;  // 219^0.35 ~= 6.594099
            8'd220: out = 12'd3382;  // 220^0.35 ~= 6.604622
            8'd221: out = 12'd3387;  // 221^0.35 ~= 6.615113
            8'd222: out = 12'd3392;  // 222^0.35 ~= 6.625574
            8'd223: out = 12'd3398;  // 223^0.35 ~= 6.636005
            8'd224: out = 12'd3403;  // 224^0.35 ~= 6.646405
            8'd225: out = 12'd3408;  // 225^0.35 ~= 6.656775
            8'd226: out = 12'd3414;  // 226^0.35 ~= 6.667115
            8'd227: out = 12'd3419;  // 227^0.35 ~= 6.677425
            8'd228: out = 12'd3424;  // 228^0.35 ~= 6.687706
            8'd229: out = 12'd3429;  // 229^0.35 ~= 6.697958
            8'd230: out = 12'd3435;  // 230^0.35 ~= 6.708181
            8'd231: out = 12'd3440;  // 231^0.35 ~= 6.718374
            8'd232: out = 12'd3445;  // 232^0.35 ~= 6.728539
            8'd233: out = 12'd3450;  // 233^0.35 ~= 6.738676
            8'd234: out = 12'd3455;  // 234^0.35 ~= 6.748784
            8'd235: out = 12'd3461;  // 235^0.35 ~= 6.758865
            8'd236: out = 12'd3466;  // 236^0.35 ~= 6.768917
            8'd237: out = 12'd3471;  // 237^0.35 ~= 6.778942
            8'd238: out = 12'd3476;  // 238^0.35 ~= 6.788939
            8'd239: out = 12'd3481;  // 239^0.35 ~= 6.798910
            8'd240: out = 12'd3486;  // 240^0.35 ~= 6.808853
            8'd241: out = 12'd3491;  // 241^0.35 ~= 6.818769
            8'd242: out = 12'd3496;  // 242^0.35 ~= 6.828658
            8'd243: out = 12'd3501;  // 243^0.35 ~= 6.838521
            8'd244: out = 12'd3506;  // 244^0.35 ~= 6.848358
            8'd245: out = 12'd3511;  // 245^0.35 ~= 6.858168
            8'd246: out = 12'd3516;  // 246^0.35 ~= 6.867953
            8'd247: out = 12'd3521;  // 247^0.35 ~= 6.877711
            8'd248: out = 12'd3526;  // 248^0.35 ~= 6.887444
            8'd249: out = 12'd3531;  // 249^0.35 ~= 6.897152
            8'd250: out = 12'd3536;  // 250^0.35 ~= 6.906834
            8'd251: out = 12'd3541;  // 251^0.35 ~= 6.916491
            8'd252: out = 12'd3546;  // 252^0.35 ~= 6.926123
            8'd253: out = 12'd3551;  // 253^0.35 ~= 6.935730
            8'd254: out = 12'd3556;  // 254^0.35 ~= 6.945313
            8'd255: out = 12'd3561;  // 255^0.35 ~= 6.954871
            default: out = 12'd0;
        endcase
    end
endmodule

// LUT for x^0.65 in Q6.6 format
module LUT_065 (
    input      [7:0] in,  // Q8.0 input
    output reg [11:0] out // Q6.6 output
);

    always @(*) begin
        case (in)
            8'd0  : out = 12'd0;  // 0^0.65 ~= 0.000000
            8'd1  : out = 12'd64;  // 1^0.65 ~= 1.000000
            8'd2  : out = 12'd100;  // 2^0.65 ~= 1.569168
            8'd3  : out = 12'd131;  // 3^0.65 ~= 2.042344
            8'd4  : out = 12'd158;  // 4^0.65 ~= 2.462289
            8'd5  : out = 12'd182;  // 5^0.65 ~= 2.846627
            8'd6  : out = 12'd205;  // 6^0.65 ~= 3.204781
            8'd7  : out = 12'd227;  // 7^0.65 ~= 3.542532
            8'd8  : out = 12'd247;  // 8^0.65 ~= 3.863745
            8'd9  : out = 12'd267;  // 9^0.65 ~= 4.171168
            8'd10 : out = 12'd286;  // 10^0.65 ~= 4.466836
            8'd11 : out = 12'd304;  // 11^0.65 ~= 4.752315
            8'd12 : out = 12'd322;  // 12^0.65 ~= 5.028840
            8'd13 : out = 12'd339;  // 13^0.65 ~= 5.297405
            8'd14 : out = 12'd356;  // 14^0.65 ~= 5.558828
            8'd15 : out = 12'd372;  // 15^0.65 ~= 5.813790
            8'd16 : out = 12'd388;  // 16^0.65 ~= 6.062866
            8'd17 : out = 12'd404;  // 17^0.65 ~= 6.306549
            8'd18 : out = 12'd419;  // 18^0.65 ~= 6.545263
            8'd19 : out = 12'd434;  // 19^0.65 ~= 6.779378
            8'd20 : out = 12'd449;  // 20^0.65 ~= 7.009217
            8'd21 : out = 12'd463;  // 21^0.65 ~= 7.235067
            8'd22 : out = 12'd477;  // 22^0.65 ~= 7.457182
            8'd23 : out = 12'd491;  // 23^0.65 ~= 7.675790
            8'd24 : out = 12'd505;  // 24^0.65 ~= 7.891096
            8'd25 : out = 12'd519;  // 25^0.65 ~= 8.103283
            8'd26 : out = 12'd532;  // 26^0.65 ~= 8.312519
            8'd27 : out = 12'd545;  // 27^0.65 ~= 8.518957
            8'd28 : out = 12'd558;  // 28^0.65 ~= 8.722736
            8'd29 : out = 12'd571;  // 29^0.65 ~= 8.923982
            8'd30 : out = 12'd584;  // 30^0.65 ~= 9.122814
            8'd31 : out = 12'd596;  // 31^0.65 ~= 9.319339
            8'd32 : out = 12'd609;  // 32^0.65 ~= 9.513657
            8'd33 : out = 12'd621;  // 33^0.65 ~= 9.705861
            8'd34 : out = 12'd633;  // 34^0.65 ~= 9.896037
            8'd35 : out = 12'd645;  // 35^0.65 ~= 10.084265
            8'd36 : out = 12'd657;  // 36^0.65 ~= 10.270619
            8'd37 : out = 12'd669;  // 37^0.65 ~= 10.455171
            8'd38 : out = 12'd681;  // 38^0.65 ~= 10.637984
            8'd39 : out = 12'd692;  // 39^0.65 ~= 10.819121
            8'd40 : out = 12'd704;  // 40^0.65 ~= 10.998640
            8'd41 : out = 12'd715;  // 41^0.65 ~= 11.176595
            8'd42 : out = 12'd727;  // 42^0.65 ~= 11.353037
            8'd43 : out = 12'd738;  // 43^0.65 ~= 11.528014
            8'd44 : out = 12'd749;  // 44^0.65 ~= 11.701573
            8'd45 : out = 12'd760;  // 45^0.65 ~= 11.873756
            8'd46 : out = 12'd771;  // 46^0.65 ~= 12.044606
            8'd47 : out = 12'd782;  // 47^0.65 ~= 12.214160
            8'd48 : out = 12'd792;  // 48^0.65 ~= 12.382456
            8'd49 : out = 12'd803;  // 49^0.65 ~= 12.549530
            8'd50 : out = 12'd814;  // 50^0.65 ~= 12.715414
            8'd51 : out = 12'd824;  // 51^0.65 ~= 12.880141
            8'd52 : out = 12'd835;  // 52^0.65 ~= 13.043741
            8'd53 : out = 12'd845;  // 53^0.65 ~= 13.206244
            8'd54 : out = 12'd856;  // 54^0.65 ~= 13.367677
            8'd55 : out = 12'd866;  // 55^0.65 ~= 13.528067
            8'd56 : out = 12'd876;  // 56^0.65 ~= 13.687440
            8'd57 : out = 12'd886;  // 57^0.65 ~= 13.845819
            8'd58 : out = 12'd896;  // 58^0.65 ~= 14.003229
            8'd59 : out = 12'd906;  // 59^0.65 ~= 14.159692
            8'd60 : out = 12'd916;  // 60^0.65 ~= 14.315229
            8'd61 : out = 12'd926;  // 61^0.65 ~= 14.469862
            8'd62 : out = 12'd936;  // 62^0.65 ~= 14.623610
            8'd63 : out = 12'd946;  // 63^0.65 ~= 14.776492
            8'd64 : out = 12'd955;  // 64^0.65 ~= 14.928528
            8'd65 : out = 12'd965;  // 65^0.65 ~= 15.079734
            8'd66 : out = 12'd975;  // 66^0.65 ~= 15.230128
            8'd67 : out = 12'd984;  // 67^0.65 ~= 15.379727
            8'd68 : out = 12'd994;  // 68^0.65 ~= 15.528546
            8'd69 : out = 12'd1003;  // 69^0.65 ~= 15.676601
            8'd70 : out = 12'd1013;  // 70^0.65 ~= 15.823907
            8'd71 : out = 12'd1022;  // 71^0.65 ~= 15.970478
            8'd72 : out = 12'd1031;  // 72^0.65 ~= 16.116329
            8'd73 : out = 12'd1041;  // 73^0.65 ~= 16.261472
            8'd74 : out = 12'd1050;  // 74^0.65 ~= 16.405921
            8'd75 : out = 12'd1059;  // 75^0.65 ~= 16.549688
            8'd76 : out = 12'd1068;  // 76^0.65 ~= 16.692786
            8'd77 : out = 12'd1077;  // 77^0.65 ~= 16.835227
            8'd78 : out = 12'd1087;  // 78^0.65 ~= 16.977021
            8'd79 : out = 12'd1096;  // 79^0.65 ~= 17.118181
            8'd80 : out = 12'd1105;  // 80^0.65 ~= 17.258716
            8'd81 : out = 12'd1114;  // 81^0.65 ~= 17.398638
            8'd82 : out = 12'd1122;  // 82^0.65 ~= 17.537957
            8'd83 : out = 12'd1131;  // 83^0.65 ~= 17.676682
            8'd84 : out = 12'd1140;  // 84^0.65 ~= 17.814824
            8'd85 : out = 12'd1149;  // 85^0.65 ~= 17.952391
            8'd86 : out = 12'd1158;  // 86^0.65 ~= 18.089393
            8'd87 : out = 12'd1166;  // 87^0.65 ~= 18.225838
            8'd88 : out = 12'd1175;  // 88^0.65 ~= 18.361736
            8'd89 : out = 12'd1184;  // 89^0.65 ~= 18.497094
            8'd90 : out = 12'd1192;  // 90^0.65 ~= 18.631921
            8'd91 : out = 12'd1201;  // 91^0.65 ~= 18.766224
            8'd92 : out = 12'd1210;  // 92^0.65 ~= 18.900012
            8'd93 : out = 12'd1218;  // 93^0.65 ~= 19.033292
            8'd94 : out = 12'd1227;  // 94^0.65 ~= 19.166072
            8'd95 : out = 12'd1235;  // 95^0.65 ~= 19.298357
            8'd96 : out = 12'd1244;  // 96^0.65 ~= 19.430157
            8'd97 : out = 12'd1252;  // 97^0.65 ~= 19.561476
            8'd98 : out = 12'd1260;  // 98^0.65 ~= 19.692323
            8'd99 : out = 12'd1269;  // 99^0.65 ~= 19.822703
            8'd100: out = 12'd1277;  // 100^0.65 ~= 19.952623
            8'd101: out = 12'd1285;  // 101^0.65 ~= 20.082089
            8'd102: out = 12'd1294;  // 102^0.65 ~= 20.211107
            8'd103: out = 12'd1302;  // 103^0.65 ~= 20.339684
            8'd104: out = 12'd1310;  // 104^0.65 ~= 20.467824
            8'd105: out = 12'd1318;  // 105^0.65 ~= 20.595533
            8'd106: out = 12'd1326;  // 106^0.65 ~= 20.722818
            8'd107: out = 12'd1334;  // 107^0.65 ~= 20.849683
            8'd108: out = 12'd1342;  // 108^0.65 ~= 20.976134
            8'd109: out = 12'd1351;  // 109^0.65 ~= 21.102175
            8'd110: out = 12'd1359;  // 110^0.65 ~= 21.227813
            8'd111: out = 12'd1367;  // 111^0.65 ~= 21.353051
            8'd112: out = 12'd1375;  // 112^0.65 ~= 21.477895
            8'd113: out = 12'd1383;  // 113^0.65 ~= 21.602350
            8'd114: out = 12'd1390;  // 114^0.65 ~= 21.726419
            8'd115: out = 12'd1398;  // 115^0.65 ~= 21.850108
            8'd116: out = 12'd1406;  // 116^0.65 ~= 21.973422
            8'd117: out = 12'd1414;  // 117^0.65 ~= 22.096364
            8'd118: out = 12'd1422;  // 118^0.65 ~= 22.218938
            8'd119: out = 12'd1430;  // 119^0.65 ~= 22.341150
            8'd120: out = 12'd1438;  // 120^0.65 ~= 22.463003
            8'd121: out = 12'd1445;  // 121^0.65 ~= 22.584501
            8'd122: out = 12'd1453;  // 122^0.65 ~= 22.705647
            8'd123: out = 12'd1461;  // 123^0.65 ~= 22.826447
            8'd124: out = 12'd1469;  // 124^0.65 ~= 22.946904
            8'd125: out = 12'd1476;  // 125^0.65 ~= 23.067021
            8'd126: out = 12'd1484;  // 126^0.65 ~= 23.186802
            8'd127: out = 12'd1492;  // 127^0.65 ~= 23.306251
            8'd128: out = 12'd1499;  // 128^0.65 ~= 23.425371
            8'd129: out = 12'd1507;  // 129^0.65 ~= 23.544166
            8'd130: out = 12'd1514;  // 130^0.65 ~= 23.662639
            8'd131: out = 12'd1522;  // 131^0.65 ~= 23.780794
            8'd132: out = 12'd1530;  // 132^0.65 ~= 23.898633
            8'd133: out = 12'd1537;  // 133^0.65 ~= 24.016160
            8'd134: out = 12'd1545;  // 134^0.65 ~= 24.133378
            8'd135: out = 12'd1552;  // 135^0.65 ~= 24.250291
            8'd136: out = 12'd1559;  // 136^0.65 ~= 24.366901
            8'd137: out = 12'd1567;  // 137^0.65 ~= 24.483211
            8'd138: out = 12'd1574;  // 138^0.65 ~= 24.599224
            8'd139: out = 12'd1582;  // 139^0.65 ~= 24.714943
            8'd140: out = 12'd1589;  // 140^0.65 ~= 24.830372
            8'd141: out = 12'd1597;  // 141^0.65 ~= 24.945512
            8'd142: out = 12'd1604;  // 142^0.65 ~= 25.060367
            8'd143: out = 12'd1611;  // 143^0.65 ~= 25.174939
            8'd144: out = 12'd1619;  // 144^0.65 ~= 25.289231
            8'd145: out = 12'd1626;  // 145^0.65 ~= 25.403245
            8'd146: out = 12'd1633;  // 146^0.65 ~= 25.516985
            8'd147: out = 12'd1640;  // 147^0.65 ~= 25.630452
            8'd148: out = 12'd1648;  // 148^0.65 ~= 25.743650
            8'd149: out = 12'd1655;  // 149^0.65 ~= 25.856580
            8'd150: out = 12'd1662;  // 150^0.65 ~= 25.969245
            8'd151: out = 12'd1669;  // 151^0.65 ~= 26.081647
            8'd152: out = 12'd1676;  // 152^0.65 ~= 26.193789
            8'd153: out = 12'd1684;  // 153^0.65 ~= 26.305674
            8'd154: out = 12'd1691;  // 154^0.65 ~= 26.417302
            8'd155: out = 12'd1698;  // 155^0.65 ~= 26.528678
            8'd156: out = 12'd1705;  // 156^0.65 ~= 26.639802
            8'd157: out = 12'd1712;  // 157^0.65 ~= 26.750677
            8'd158: out = 12'd1719;  // 158^0.65 ~= 26.861305
            8'd159: out = 12'd1726;  // 159^0.65 ~= 26.971688
            8'd160: out = 12'd1733;  // 160^0.65 ~= 27.081829
            8'd161: out = 12'd1740;  // 161^0.65 ~= 27.191729
            8'd162: out = 12'd1747;  // 162^0.65 ~= 27.301390
            8'd163: out = 12'd1754;  // 163^0.65 ~= 27.410815
            8'd164: out = 12'd1761;  // 164^0.65 ~= 27.520005
            8'd165: out = 12'd1768;  // 165^0.65 ~= 27.628962
            8'd166: out = 12'd1775;  // 166^0.65 ~= 27.737688
            8'd167: out = 12'd1782;  // 167^0.65 ~= 27.846185
            8'd168: out = 12'd1789;  // 168^0.65 ~= 27.954455
            8'd169: out = 12'd1796;  // 169^0.65 ~= 28.062500
            8'd170: out = 12'd1803;  // 170^0.65 ~= 28.170321
            8'd171: out = 12'd1810;  // 171^0.65 ~= 28.277921
            8'd172: out = 12'd1817;  // 172^0.65 ~= 28.385300
            8'd173: out = 12'd1824;  // 173^0.65 ~= 28.492461
            8'd174: out = 12'd1830;  // 174^0.65 ~= 28.599406
            8'd175: out = 12'd1837;  // 175^0.65 ~= 28.706136
            8'd176: out = 12'd1844;  // 176^0.65 ~= 28.812652
            8'd177: out = 12'd1851;  // 177^0.65 ~= 28.918957
            8'd178: out = 12'd1858;  // 178^0.65 ~= 29.025052
            8'd179: out = 12'd1864;  // 179^0.65 ~= 29.130938
            8'd180: out = 12'd1871;  // 180^0.65 ~= 29.236618
            8'd181: out = 12'd1878;  // 181^0.65 ~= 29.342092
            8'd182: out = 12'd1885;  // 182^0.65 ~= 29.447362
            8'd183: out = 12'd1891;  // 183^0.65 ~= 29.552431
            8'd184: out = 12'd1898;  // 184^0.65 ~= 29.657298
            8'd185: out = 12'd1905;  // 185^0.65 ~= 29.761966
            8'd186: out = 12'd1911;  // 186^0.65 ~= 29.866437
            8'd187: out = 12'd1918;  // 187^0.65 ~= 29.970711
            8'd188: out = 12'd1925;  // 188^0.65 ~= 30.074790
            8'd189: out = 12'd1931;  // 189^0.65 ~= 30.178675
            8'd190: out = 12'd1938;  // 190^0.65 ~= 30.282369
            8'd191: out = 12'd1945;  // 191^0.65 ~= 30.385871
            8'd192: out = 12'd1951;  // 192^0.65 ~= 30.489184
            8'd193: out = 12'd1958;  // 193^0.65 ~= 30.592309
            8'd194: out = 12'd1964;  // 194^0.65 ~= 30.695246
            8'd195: out = 12'd1971;  // 195^0.65 ~= 30.797999
            8'd196: out = 12'd1978;  // 196^0.65 ~= 30.900567
            8'd197: out = 12'd1984;  // 197^0.65 ~= 31.002952
            8'd198: out = 12'd1991;  // 198^0.65 ~= 31.105155
            8'd199: out = 12'd1997;  // 199^0.65 ~= 31.207178
            8'd200: out = 12'd2004;  // 200^0.65 ~= 31.309022
            8'd201: out = 12'd2010;  // 201^0.65 ~= 31.410687
            8'd202: out = 12'd2017;  // 202^0.65 ~= 31.512176
            8'd203: out = 12'd2023;  // 203^0.65 ~= 31.613489
            8'd204: out = 12'd2030;  // 204^0.65 ~= 31.714627
            8'd205: out = 12'd2036;  // 205^0.65 ~= 31.815592
            8'd206: out = 12'd2043;  // 206^0.65 ~= 31.916385
            8'd207: out = 12'd2049;  // 207^0.65 ~= 32.017007
            8'd208: out = 12'd2056;  // 208^0.65 ~= 32.117458
            8'd209: out = 12'd2062;  // 209^0.65 ~= 32.217741
            8'd210: out = 12'd2068;  // 210^0.65 ~= 32.317856
            8'd211: out = 12'd2075;  // 211^0.65 ~= 32.417804
            8'd212: out = 12'd2081;  // 212^0.65 ~= 32.517587
            8'd213: out = 12'd2088;  // 213^0.65 ~= 32.617205
            8'd214: out = 12'd2094;  // 214^0.65 ~= 32.716659
            8'd215: out = 12'd2100;  // 215^0.65 ~= 32.815951
            8'd216: out = 12'd2107;  // 216^0.65 ~= 32.915082
            8'd217: out = 12'd2113;  // 217^0.65 ~= 33.014052
            8'd218: out = 12'd2119;  // 218^0.65 ~= 33.112862
            8'd219: out = 12'd2126;  // 219^0.65 ~= 33.211514
            8'd220: out = 12'd2132;  // 220^0.65 ~= 33.310008
            8'd221: out = 12'd2138;  // 221^0.65 ~= 33.408346
            8'd222: out = 12'd2144;  // 222^0.65 ~= 33.506528
            8'd223: out = 12'd2151;  // 223^0.65 ~= 33.604556
            8'd224: out = 12'd2157;  // 224^0.65 ~= 33.702430
            8'd225: out = 12'd2163;  // 225^0.65 ~= 33.800151
            8'd226: out = 12'd2169;  // 226^0.65 ~= 33.897720
            8'd227: out = 12'd2176;  // 227^0.65 ~= 33.995138
            8'd228: out = 12'd2182;  // 228^0.65 ~= 34.092406
            8'd229: out = 12'd2188;  // 229^0.65 ~= 34.189525
            8'd230: out = 12'd2194;  // 230^0.65 ~= 34.286495
            8'd231: out = 12'd2201;  // 231^0.65 ~= 34.383318
            8'd232: out = 12'd2207;  // 232^0.65 ~= 34.479995
            8'd233: out = 12'd2213;  // 233^0.65 ~= 34.576525
            8'd234: out = 12'd2219;  // 234^0.65 ~= 34.672911
            8'd235: out = 12'd2225;  // 235^0.65 ~= 34.769153
            8'd236: out = 12'd2231;  // 236^0.65 ~= 34.865251
            8'd237: out = 12'd2238;  // 237^0.65 ~= 34.961208
            8'd238: out = 12'd2244;  // 238^0.65 ~= 35.057022
            8'd239: out = 12'd2250;  // 239^0.65 ~= 35.152696
            8'd240: out = 12'd2256;  // 240^0.65 ~= 35.248229
            8'd241: out = 12'd2262;  // 241^0.65 ~= 35.343624
            8'd242: out = 12'd2268;  // 242^0.65 ~= 35.438880
            8'd243: out = 12'd2274;  // 243^0.65 ~= 35.533998
            8'd244: out = 12'd2280;  // 244^0.65 ~= 35.628980
            8'd245: out = 12'd2286;  // 245^0.65 ~= 35.723825
            8'd246: out = 12'd2292;  // 246^0.65 ~= 35.818535
            8'd247: out = 12'd2298;  // 247^0.65 ~= 35.913110
            8'd248: out = 12'd2304;  // 248^0.65 ~= 36.007552
            8'd249: out = 12'd2311;  // 249^0.65 ~= 36.101860
            8'd250: out = 12'd2317;  // 250^0.65 ~= 36.196036
            8'd251: out = 12'd2323;  // 251^0.65 ~= 36.290079
            8'd252: out = 12'd2329;  // 252^0.65 ~= 36.383992
            8'd253: out = 12'd2335;  // 253^0.65 ~= 36.477775
            8'd254: out = 12'd2341;  // 254^0.65 ~= 36.571428
            8'd255: out = 12'd2347;  // 255^0.65 ~= 36.664952
            default: out = 12'd0;
        endcase
    end
endmodule
